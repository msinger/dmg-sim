`default_nettype none

module sm83_nor2_in2_n #(
		parameter real L_y = 8
	) (
		input  logic in1, in2_n,
		output logic y
	);

	import sm83_timing::*;

	assign y = !(in1 | !in2_n);

	specify
		specparam T_rise_in2 = tpd_elmore( 28, R_pmos_ohm(3*L_unit));
		specparam T_fall_in2 = tpd_elmore( 28, R_nmos_ohm(3*L_unit));
		specparam T_rise_y   = tpd_elmore(L_y, R_pmos_ohm(3*L_unit) * 2);
		specparam T_fall_y   = tpd_elmore(L_y, R_nmos_ohm(3*L_unit));

		(in1   *> y) = (T_rise_y, T_fall_y);
		(in2_n *> y) = (T_fall_in2 + T_rise_y, T_rise_in2 + T_fall_y);
	endspecify

endmodule

`default_nettype wire
