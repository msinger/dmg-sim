`default_nettype none

module sprite_x_matchers(
		inout tri logic [7:0] d,
		input logic     [7:0] oam_a_nd, nh,

		input logic clk3, oam_a_cpu_nrd,
		input logic cota, dyna, fuxu, wupa, yfag, gafy, gecy, asys, doku, zape, xaho, wunu, wofo,
		input logic wuzo, cexu, dosy, weme, ejad, cyla, cacu, gamy,

		output logic ngomo, nbaxo, nyzos, ndepo, xeba, zako, ywos, zure, daje, cyco, cyvy, ewam,
		output logic ywap, ydot, ykok, ynaz, dama, feha, ytub, ylev, cogy, fyma, cehu, ekes
	);

	logic wyno, cyra, zuve, eced, xyky, yrum, ysex, yvel;
	logic xega, gomo, baxo, yzos, depo, ylor, zyty, zyve, zezy;
	logic cose, arop, xatu, bady, zago, zocy, ypur, yvok;
	logic xaca, xagu, xepu, xygu, xuna, deve, zeha, fyra;
	logic welo, xuny, wote, xako, xepe, ylah, zola, zulu;
	logic woju, yfun, wyza, ypuk, zogy, zeba, zaha, zoky;
	logic xomy, wuha, wyna, weco, xoly, xyba, xabe, xeka;
	logic yvap, xeny, xavu, xeva, yhok, ycah, ydaj, yvuz;
	logic fazu, faxe, exuk, fede, eraz, epum, erol, ehyn;
	logic ejot, esaj, ducu, ewud, duse, dagu, dyze, deso;
	logic dake, ceso, dyfu, cusy, dany, duko, desu, dazo;
	logic cola, boba, colu, bahu, edym, emyb, ebef, ewok;
	logic zoly, zogo, zecu, zesa, ycol, yrac, ymem, yvag;
	logic zare, zemu, zygo, zuzy, xosu, zuvu, xuco, zulo;
	logic ybed, zala, wyde, xepa, wedu, ygaj, zyjo, xury;
	logic zyku, zypu, xaha, zefe, xeju, zate, zaku, ybox;
	logic ezuf, enad, ebow, fyca, gavy, gypu, gady, gaza;
	logic duze, daga, dawu, ejaw, goho, gasu, gabu, gafe;
	logic ypod, yrop, ynep, yzof, xuvy, xere, xuzo, xexa;
	logic zywu, zuza, zejo, zeda, ymam, ytyp, yfop, yvac;
	logic cywe, dyby, dury, cuvy, fusa, faxa, fozy, fesy;
	logic bazy, cyle, ceva, bumy, guzo, gola, geve, gude;
	logic duhy, ejuf, enor, depy, foka, fyty, fuby, goxu;
	logic ceko, dety, dozo, cony, fuzu, feso, foky, fyva;
	dlatch latch_wyno(clk3, oam_a_nd[4], wyno);
	dlatch latch_cyra(clk3, oam_a_nd[5], cyra);
	dlatch latch_zuve(clk3, oam_a_nd[6], zuve);
	dlatch latch_eced(clk3, oam_a_nd[7], eced);
	dlatch latch_xyky(clk3, oam_a_nd[0], xyky);
	dlatch latch_yrum(clk3, oam_a_nd[1], yrum);
	dlatch latch_ysex(clk3, oam_a_nd[2], ysex);
	dlatch latch_yvel(clk3, oam_a_nd[3], yvel);
	dff dff_gomo(xega, wyno, gomo);
	dff dff_baxo(xega, cyra, baxo);
	dff dff_yzos(xega, zuve, yzos);
	dff dff_depo(xega, eced, depo);
	dff dff_ylor(xega, xyky, ylor);
	dff dff_zyty(xega, yrum, zyty);
	dff dff_zyve(xega, ysex, zyve);
	dff dff_zezy(xega, yvel, zezy);
	dffr_a dffr_welo(fuxu, dyna, cose, welo);
	dffr_a dffr_xuny(fuxu, dyna, arop, xuny);
	dffr_a dffr_wote(fuxu, dyna, xatu, wote);
	dffr_a dffr_xako(fuxu, dyna, bady, xako);
	dffr_a dffr_xepe(fuxu, dyna, zago, xepe);
	dffr_a dffr_ylah(fuxu, dyna, zocy, ylah);
	dffr_a dffr_zola(fuxu, dyna, ypur, zola);
	dffr_a dffr_zulu(fuxu, dyna, yvok, zulu);
	dffr_a dffr_xomy(yfag, wupa, cose, xomy);
	dffr_a dffr_wuha(yfag, wupa, arop, wuha);
	dffr_a dffr_wyna(yfag, wupa, xatu, wyna);
	dffr_a dffr_weco(yfag, wupa, bady, weco);
	dffr_a dffr_xoly(yfag, wupa, zago, xoly);
	dffr_a dffr_xyba(yfag, wupa, zocy, xyba);
	dffr_a dffr_xabe(yfag, wupa, ypur, xabe);
	dffr_a dffr_xeka(yfag, wupa, yvok, xeka);
	dffr_a dffr_fazu(gecy, gafy, cose, fazu);
	dffr_a dffr_faxe(gecy, gafy, arop, faxe);
	dffr_a dffr_exuk(gecy, gafy, xatu, exuk);
	dffr_a dffr_fede(gecy, gafy, bady, fede);
	dffr_a dffr_eraz(gecy, gafy, zago, eraz);
	dffr_a dffr_epum(gecy, gafy, zocy, epum);
	dffr_a dffr_erol(gecy, gafy, ypur, erol);
	dffr_a dffr_ehyn(gecy, gafy, yvok, ehyn);
	dffr_a dffr_dake(asys, doku, cose, dake);
	dffr_a dffr_ceso(asys, doku, arop, ceso);
	dffr_a dffr_dyfu(asys, doku, xatu, dyfu);
	dffr_a dffr_cusy(asys, doku, bady, cusy);
	dffr_a dffr_dany(asys, doku, zago, dany);
	dffr_a dffr_duko(asys, doku, zocy, duko);
	dffr_a dffr_desu(asys, doku, ypur, desu);
	dffr_a dffr_dazo(asys, doku, yvok, dazo);
	dffr_a dffr_zoly(zape, xaho, cose, zoly);
	dffr_a dffr_zogo(zape, xaho, arop, zogo);
	dffr_a dffr_zecu(zape, xaho, xatu, zecu);
	dffr_a dffr_zesa(zape, xaho, bady, zesa);
	dffr_a dffr_ycol(zape, xaho, zago, ycol);
	dffr_a dffr_yrac(zape, xaho, zocy, yrac);
	dffr_a dffr_ymem(zape, xaho, ypur, ymem);
	dffr_a dffr_yvag(zape, xaho, yvok, yvag);
	dffr_a dffr_ybed(wofo, wunu, cose, ybed);
	dffr_a dffr_zala(wofo, wunu, arop, zala);
	dffr_a dffr_wyde(wofo, wunu, xatu, wyde);
	dffr_a dffr_xepa(wofo, wunu, bady, xepa);
	dffr_a dffr_wedu(wofo, wunu, zago, wedu);
	dffr_a dffr_ygaj(wofo, wunu, zocy, ygaj);
	dffr_a dffr_zyjo(wofo, wunu, ypur, zyjo);
	dffr_a dffr_xury(wofo, wunu, yvok, xury);
	dffr_a dffr_ezuf(cexu, wuzo, cose, ezuf);
	dffr_a dffr_enad(cexu, wuzo, arop, enad);
	dffr_a dffr_ebow(cexu, wuzo, xatu, ebow);
	dffr_a dffr_fyca(cexu, wuzo, bady, fyca);
	dffr_a dffr_gavy(cexu, wuzo, zago, gavy);
	dffr_a dffr_gypu(cexu, wuzo, zocy, gypu);
	dffr_a dffr_gady(cexu, wuzo, ypur, gady);
	dffr_a dffr_gaza(cexu, wuzo, yvok, gaza);
	dffr_a dffr_ypod(weme, dosy, cose, ypod);
	dffr_a dffr_yrop(weme, dosy, arop, yrop);
	dffr_a dffr_ynep(weme, dosy, xatu, ynep);
	dffr_a dffr_yzof(weme, dosy, bady, yzof);
	dffr_a dffr_xuvy(weme, dosy, zago, xuvy);
	dffr_a dffr_xere(weme, dosy, zocy, xere);
	dffr_a dffr_xuzo(weme, dosy, ypur, xuzo);
	dffr_a dffr_xexa(weme, dosy, yvok, xexa);
	dffr_a dffr_cywe(cyla, ejad, cose, cywe);
	dffr_a dffr_dyby(cyla, ejad, arop, dyby);
	dffr_a dffr_dury(cyla, ejad, xatu, dury);
	dffr_a dffr_cuvy(cyla, ejad, bady, cuvy);
	dffr_a dffr_fusa(cyla, ejad, zago, fusa);
	dffr_a dffr_faxa(cyla, ejad, zocy, faxa);
	dffr_a dffr_fozy(cyla, ejad, ypur, fozy);
	dffr_a dffr_fesy(cyla, ejad, yvok, fesy);
	dffr_a dffr_duhy(cacu, gamy, cose, duhy);
	dffr_a dffr_ejuf(cacu, gamy, arop, ejuf);
	dffr_a dffr_enor(cacu, gamy, xatu, enor);
	dffr_a dffr_depy(cacu, gamy, bady, depy);
	dffr_a dffr_foka(cacu, gamy, zago, foka);
	dffr_a dffr_fyty(cacu, gamy, zocy, fyty);
	dffr_a dffr_fuby(cacu, gamy, ypur, fuby);
	dffr_a dffr_goxu(cacu, gamy, yvok, goxu);
	assign #T_INV  xega = !cota;
	assign #T_INV  cose = !(!gomo);
	assign #T_INV  arop = !(!baxo);
	assign #T_INV  xatu = !(!yzos);
	assign #T_INV  bady = !(!depo);
	assign #T_INV  zago = !(!ylor);
	assign #T_INV  zocy = !(!zyty);
	assign #T_INV  ypur = !(!zyve);
	assign #T_INV  yvok = !(!zezy);
	assign #T_TRIB xaca = !oam_a_cpu_nrd ? !xyky : 'z;
	assign #T_TRIB xagu = !oam_a_cpu_nrd ? !yrum : 'z;
	assign #T_TRIB xepu = !oam_a_cpu_nrd ? !ysex : 'z;
	assign #T_TRIB xygu = !oam_a_cpu_nrd ? !yvel : 'z;
	assign #T_TRIB xuna = !oam_a_cpu_nrd ? !wyno : 'z;
	assign #T_TRIB deve = !oam_a_cpu_nrd ? !cyra : 'z;
	assign #T_TRIB zeha = !oam_a_cpu_nrd ? !zuve : 'z;
	assign #T_TRIB fyra = !oam_a_cpu_nrd ? !eced : 'z;
	assign #T_XOR  woju = welo != nh[4];
	assign #T_XOR  yfun = xuny != nh[5];
	assign #T_XOR  wyza = wote != nh[6];
	assign #T_XOR  ypuk = xako != nh[7];
	assign #T_XOR  zogy = xepe != nh[0];
	assign #T_XOR  zeba = ylah != nh[1];
	assign #T_XOR  zaha = zola != nh[2];
	assign #T_XOR  zoky = zulu != nh[3];
	assign #T_NOR  xeba = !(woju || yfun || wyza || ypuk);
	assign #T_NOR  zako = !(zogy || zeba || zaha || zoky);
	assign #T_XOR  yvap = xomy != nh[4];
	assign #T_XOR  xeny = wuha != nh[5];
	assign #T_XOR  xavu = wyna != nh[6];
	assign #T_XOR  xeva = weco != nh[7];
	assign #T_XOR  yhok = xoly != nh[0];
	assign #T_XOR  ycah = xyba != nh[1];
	assign #T_XOR  ydaj = xabe != nh[2];
	assign #T_XOR  yvuz = xeka != nh[3];
	assign #T_NOR  ywos = !(yvap || xeny || xavu || xeva);
	assign #T_NOR  zure = !(yhok || ycah || ydaj || yvuz);
	assign #T_XOR  ejot = fazu != nh[4];
	assign #T_XOR  esaj = faxe != nh[5];
	assign #T_XOR  ducu = exuk != nh[6];
	assign #T_XOR  ewud = fede != nh[7];
	assign #T_XOR  duse = eraz != nh[0];
	assign #T_XOR  dagu = epum != nh[1];
	assign #T_XOR  dyze = erol != nh[2];
	assign #T_XOR  deso = ehyn != nh[3];
	assign #T_NOR  daje = !(ejot || esaj || ducu || ewud);
	assign #T_NOR  cyco = !(duse || dagu || dyze || deso);
	assign #T_XOR  cola = dake != nh[4];
	assign #T_XOR  boba = ceso != nh[5];
	assign #T_XOR  colu = dyfu != nh[6];
	assign #T_XOR  bahu = cusy != nh[7];
	assign #T_XOR  edym = dany != nh[0];
	assign #T_XOR  emyb = duko != nh[1];
	assign #T_XOR  ebef = desu != nh[2];
	assign #T_XOR  ewok = dazo != nh[3];
	assign #T_NOR  cyvy = !(cola || boba || colu || bahu);
	assign #T_NOR  ewam = !(edym || emyb || ebef || ewok);
	assign #T_XOR  zare = zoly != nh[4];
	assign #T_XOR  zemu = zogo != nh[5];
	assign #T_XOR  zygo = zecu != nh[6];
	assign #T_XOR  zuzy = zesa != nh[7];
	assign #T_XOR  xosu = ycol != nh[0];
	assign #T_XOR  zuvu = yrac != nh[1];
	assign #T_XOR  xuco = ymem != nh[2];
	assign #T_XOR  zulo = yvag != nh[3];
	assign #T_NOR  ywap = !(zare || zemu || zygo || zuzy);
	assign #T_NOR  ydot = !(xosu || zuvu || xuco || zulo);
	assign #T_XOR  zyku = ybed != nh[4];
	assign #T_XOR  zypu = zala != nh[5];
	assign #T_XOR  xaha = wyde != nh[6];
	assign #T_XOR  zefe = xepa != nh[7];
	assign #T_XOR  xeju = wedu != nh[0];
	assign #T_XOR  zate = ygaj != nh[1];
	assign #T_XOR  zaku = zyjo != nh[2];
	assign #T_XOR  ybox = xury != nh[3];
	assign #T_NOR  ykok = !(zyku || zypu || xaha || zefe);
	assign #T_NOR  ynaz = !(xeju || zate || zaku || ybox);
	assign #T_XOR  duze = ezuf != nh[4];
	assign #T_XOR  daga = enad != nh[5];
	assign #T_XOR  dawu = ebow != nh[6];
	assign #T_XOR  ejaw = fyca != nh[7];
	assign #T_XOR  goho = gavy != nh[0];
	assign #T_XOR  gasu = gypu != nh[1];
	assign #T_XOR  gabu = gady != nh[2];
	assign #T_XOR  gafe = gaza != nh[3];
	assign #T_NOR  dama = !(duze || daga || dawu || ejaw);
	assign #T_NOR  feha = !(goho || gasu || gabu || gafe);
	assign #T_XOR  zywu = ypod != nh[4];
	assign #T_XOR  zuza = yrop != nh[5];
	assign #T_XOR  zejo = ynep != nh[6];
	assign #T_XOR  zeda = yzof != nh[7];
	assign #T_XOR  ymam = xuvy != nh[0];
	assign #T_XOR  ytyp = xere != nh[1];
	assign #T_XOR  yfop = xuzo != nh[2];
	assign #T_XOR  yvac = xexa != nh[3];
	assign #T_NOR  ytub = !(zywu || zuza || zejo || zeda);
	assign #T_NOR  ylev = !(ymam || ytyp || yfop || yvac);
	assign #T_XOR  bazy = cywe != nh[4];
	assign #T_XOR  cyle = dyby != nh[5];
	assign #T_XOR  ceva = dury != nh[6];
	assign #T_XOR  bumy = cuvy != nh[7];
	assign #T_XOR  guzo = fusa != nh[0];
	assign #T_XOR  gola = faxa != nh[1];
	assign #T_XOR  geve = fozy != nh[2];
	assign #T_XOR  gude = fesy != nh[3];
	assign #T_NOR  cogy = !(bazy || cyle || ceva || bumy);
	assign #T_NOR  fyma = !(guzo || gola || geve || gude);
	assign #T_XOR  ceko = duhy != nh[4];
	assign #T_XOR  dety = ejuf != nh[5];
	assign #T_XOR  dozo = enor != nh[6];
	assign #T_XOR  cony = depy != nh[7];
	assign #T_XOR  fuzu = foka != nh[0];
	assign #T_XOR  feso = fyty != nh[1];
	assign #T_XOR  foky = fuby != nh[2];
	assign #T_XOR  fyva = goxu != nh[3];
	assign #T_NOR  cehu = !(ceko || dety || dozo || cony);
	assign #T_NOR  ekes = !(fuzu || feso || foky || fyva);
	assign ngomo = !gomo;
	assign nbaxo = !baxo;
	assign nyzos = !yzos;
	assign ndepo = !depo;
	assign d[0] = xaca;
	assign d[1] = xagu;
	assign d[2] = xepu;
	assign d[3] = xygu;
	assign d[4] = xuna;
	assign d[5] = deve;
	assign d[6] = zeha;
	assign d[7] = fyra;

endmodule
