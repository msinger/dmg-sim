`default_nettype none
`timescale 1ns/100ps

parameter T_INV   = 2;
parameter T_AND   = 4;
parameter T_NAND  = 2;
parameter T_OR    = 4;
parameter T_NOR   = 2;
parameter T_OA    = 6;
parameter T_AO    = 6;
parameter T_NAO   = 5;
parameter T_MUX   = 6;
parameter T_TRI   = 2;
parameter T_DFFR  = 8;
parameter T_DFF   = 8;
parameter T_LATCH = 4;

module dmg;

	reg [31:0] cyc;

	reg xi;
	wire clkin_a, clkin_b;
	wire reset; /* inverted !RST pin */
	wire t1 = 0;
	wire t2 = 0;
	assign clkin_a = cyc >= 2;
	assign clkin_b = xi;
	assign reset = cyc >= 40 && cyc <= 80;

	initial begin
		$dumpfile("dmg.vcd");
		$dumpvars(0, dmg);

		cyc = 0;
		xi  = 0;
	end

	always #122 xi = !xi;

	always @(posedge xi) begin
		cyc++;
		if (cyc == 10000) $finish;
	end

	wire [7:0]  d, d_a, d_d, md, md_out, md_a, oam_a_d, oam_b_d;
	wire [15:0] a, a_a, a_d, dma_a;
	wire [12:0] ma, ma_out;

	wire wr_a, wr_c, rd_a, rd_c;
	wire moe_a, moe_d, mwr_a, mwr_d, mcs_a, mcs_d, md_b;

	assign a = 0;

	/* not yet generated signals */
	wire [7:0] d_in = 'hff;
	wire [7:0] md_in = 'hff;
	wire [15:0] a_c = 0;
	wire wr_in = 0;
	wire rd_b = 0;
	wire moe_in = 0;
	wire mwr_in = 0;
	wire mcs_in = 0;
	wire cpu_raw_rd = 0;
	wire cpu_wr_raw = 0;
	wire ff40_d7 = 0;
	wire from_cpu = 0;
	wire from_cpu3 = 1;
	wire from_cpu4 = 0;
	wire from_cpu5 = 0;
	wire from_cpu6 = 0;
	wire clk_from_cpu = 1;
	wire tovy_na0 = 1;
	wire a00_07 = 0;
	wire ff46 = 0;
	wire ff40_d4 = 0;
	wire amab = 0;
	wire nff1a_d7 = 1;
	wire nch1_amp_en = 1;
	wire nch2_amp_en = 1;
	wire nch4_amp_en = 1;
	wire nch1_active = 1;
	wire nch2_active = 1;
	wire nch3_active = 1;
	wire nch4_active = 1;
	wire tacu = 0;
	wire tuvo = 0;
	wire acyl = 0;
	wire xyso = 0;
	wire texy = 0;
	wire myma = 0;
	wire lena = 0;
	wire xymu = 0;
	wire leko = 0;
	wire xuha = 0;
	wire vyno = 0;
	wire vujo = 0;
	wire vymu = 0;
	wire neta = 0;
	wire pore = 0;
	wire potu = 0;
	wire npyju = 1;
	wire npowy = 1;
	wire npoju = 1;
	wire npulo = 1;
	wire npoxa = 1;
	wire npyzo = 1;
	wire npozo = 1;
	wire nrawu = 1;

	wire clk1;

	wire cpu_wr, cpu_wr2;
	wire cpu_rd, cpu_rd2;
	wire cpu_rd_sync;
	wire nt1_nt2, nt1_t2, t1_nt2;
	wire ff04_ff07, ff0f_rd, ff0f_wr, ff00wr, ff00rd;
	wire apu_wr, ncpu_rd;
	wire hram_cs, boot_cs, ncs_out;
	wire to_cpu, to_cpu_tutu;

	wire nreset2, nreset6;
	wire nphi_out;

	wire dma_run, vram_to_oam, dma_addr_ext, oam_addr_dma;
	wire caty, wyja, mopa_phi;
	wire tola_na1;

	wire ff60_d1, ff60_d0;
	wire ff26, ff3x, namp_en;

	wire apu_reset, net03;
	wire napu_reset, napu_reset2, napu_reset4, napu_reset5, napu_reset6;
	wire apuv_4mhz;
	wire ajer_2mhz;
	wire byfe_128hz;
	wire dyfa_1mhz;
	wire afas, fero_q, cate, gaxo, bedo, abuz, tutu, texo, roru, lula, anap, duce, cota, wuko;

	wire ffxx, nffxx, nfexxffxx, saro;
	wire ff10, ff11, ff12, ff13, ff14, ff16, ff17, ff18, ff19, ff1a;
	wire ff1b, ff1c, ff1d, ff1e, ff20, ff21, ff22, ff23, ff24, ff25;

	wire [3:0] lmixer, rmixer;

	clk            p1_clk(.*);
	dma            p4_dma(.*);
	sys_decode     p7_sys_decode(.*);
	ext_cpu_busses p8_ext_cpu_busses(.*);
	apu_ctrl       p9_apu_ctrl(.*);
	apu_decode     p10_apu_decode(.*);
	vram_ifc       p25_vram_ifc(.*);

endmodule

module clk(
		clkin_a, clkin_b, reset,
		nreset2, nreset6,
		clk1, nphi_out,
		d,
		cpu_rd_sync,
		cpu_wr, cpu_rd,
		nt1_nt2, nt1_t2, t1_nt2,
		from_cpu3, from_cpu4, clk_from_cpu, to_cpu,
		ff04_ff07, ff40_d7, ff60_d1, tovy_na0, tola_na1,
		apu_reset, napu_reset5,
		apuv_4mhz, ajer_2mhz, byfe_128hz,
		fero_q, bedo, abuz, afas
	);

	input wire clkin_a, clkin_b;
	input wire reset;

	output wire nreset2, nreset6;
	output wire clk1;
	output wire nphi_out;

	inout wire [7:0] d;

	output wire cpu_rd_sync;
	input  wire cpu_wr, cpu_rd;
	input  wire nt1_nt2, nt1_t2, t1_nt2;

	input  wire from_cpu3;
	input  wire from_cpu4;
	input  wire clk_from_cpu;
	output wire to_cpu;

	input wire ff04_ff07;
	input wire ff40_d7;
	input wire ff60_d1;
	input wire tovy_na0;
	input wire tola_na1;

	input  wire apu_reset;
	input  wire napu_reset5;
	output wire apuv_4mhz;
	input  wire ajer_2mhz;
	output wire byfe_128hz;
	input  wire fero_q;
	output wire bedo, abuz, afas;

	wire arys, anos, avet;
	assign #T_INV  arys = !clkin_b;
	assign #T_NAND anos = !(clkin_b && avet);
	assign #T_NAND avet = !(anos && arys);

	wire atal, atal_4mhz;
	assign #T_INV  atal = !avet;
	assign atal_4mhz = atal;

	wire azof, zaxy, zeme, alet, lape, tava, atag, amuk, clk2, clk4, clk5, amuk_4mhz;
	assign #T_INV  azof = !atal;
	assign #T_INV  zaxy = !azof;
	assign #T_INV  zeme = !zaxy;
	assign #T_INV  alet = !zeme;
	assign #T_INV  lape = !alet;
	assign #T_INV  tava = !lape;
	assign #T_INV  atag = !azof;
	assign #T_INV  amuk = !atag;
	assign clk1 = zeme;
	assign clk2 = alet;
	assign clk4 = lape;
	assign clk5 = tava;
	assign amuk_4mhz = amuk;

	wire aryf, apuv, cybo, bela, cery, aryf_4mhz, cery_2mhz;
	assign #T_INV  aryf = !amuk;
	assign #T_INV  apuv = !amuk;
	assign #T_INV  cybo = !amuk;
	assign #T_INV  bela = !apu_reset;
	dffr dffr_cery(cybo, bela, !cery, cery);
	assign aryf_4mhz = aryf;
	assign apuv_4mhz = apuv;
	assign cery_2mhz = cery;

	wire dula, cunu, xore, walu, wesy, xebe, reset7, nreset7, nreset8, nreset9;
	assign #T_INV  dula = !nreset2;
	assign #T_INV  cunu = !dula;
	assign #T_INV  xore = !cunu;
	assign #T_INV  walu = !xore;
	assign #T_INV  wesy = !xore;
	assign #T_INV  xebe = !xore;
	assign nreset6 = cunu;
	assign reset7  = xore;
	assign nreset7 = xebe;
	assign nreset8 = walu;
	assign nreset9 = wesy;

	wire xodo, xapo, pyry, atar, lyha, lyfe, reset_video, nreset_video, reset_video2, nreset_video2, reset_video3;
	assign #T_NAND xodo = !(ff40_d7 && nreset7);
	assign #T_INV  xapo = !xodo;
	assign #T_INV  pyry = !xapo;
	assign #T_INV  atar = !xapo;
	assign #T_INV  lyha = !xapo;
	assign #T_INV  lyfe = !lyha;
	assign reset_video   = atar;
	assign nreset_video  = xapo;
	assign reset_video2  = pyry;
	assign nreset_video2 = lyfe;
	assign reset_video3  = lyha;

	wire adyk, afur, alef, apuk, abol, ucob, uvyt, nclkin_a;
	wire adar, atyp, afep, arov, ajax, bugo, arev, apov, agut, awod, bate, basu, buke;
	dffr dffr_adyk(atal_4mhz,  nt1_nt2, apuk,  adyk);
	dffr dffr_afur(!atal_4mhz, nt1_nt2, !adyk, afur);
	dffr dffr_alef(atal_4mhz,  nt1_nt2, afur,  alef);
	dffr dffr_apuk(!atal_4mhz, nt1_nt2, alef,  apuk);
	assign #T_INV  abol = !clk_from_cpu;
	assign #T_INV  ucob = !clkin_a;
	assign #T_INV  uvyt = !phi_out;
	assign #T_INV  adar = !adyk;
	assign #T_INV  atyp = afur; /* takes !q output of dff */
	assign #T_INV  afep = !alef;
	assign #T_INV  arov = apuk; /* takes !q output of dff */
	assign #T_NOR  afas = !(adar || atyp);
	assign #T_NAND arev = !(from_cpu3 && afas);
	assign #T_INV  apov = !arev;
	assign #T_INV  ajax = !atyp;
	assign #T_INV  bugo = !afep;
	assign #T_OA   agut = (ajax || arov) && from_cpu4;
	assign #T_OR   awod = nt1_t2 || agut;
	assign #T_INV  abuz = !awod;
	assign #T_NOR  bate = !(bugo || arov || abol);
	assign #T_INV  basu = !bate;
	assign #T_INV  buke = !basu;
	assign nclkin_a = ucob;
	assign nphi_out = uvyt;
	assign cpu_rd_sync = apov;

	wire bapy, belu, beru, byry, bufa, byly, bude, beva, bolo, byda, beko, bavy, beja, dova, phi_out, nphi;
	wire bane, belo, baze, buto;
	assign #T_NOR  bapy = !(abol || arov || atyp);
	assign #T_NOR  belu = !(atyp || abol);
	assign #T_INV  beru = !bapy;
	assign #T_INV  byry = !belu;
	assign #T_INV  bufa = !beru;
	assign #T_INV  byly = !beru;
	assign #T_INV  bude = !byry;
	assign #T_INV  beva = !byry;
	assign #T_INV  bolo = !bufa;
	assign #T_INV  byda = !bufa;
	assign #T_INV  beko = !bude;
	assign #T_INV  bavy = !bude;
	assign #T_INV  dova = !bude;
	assign #T_NAND beja = !(bolo && beko);
	assign #T_INV  bane = !beja;
	assign #T_INV  belo = !bane;
	assign #T_INV  baze = !belo;
	assign #T_NAND buto = !(afep && atyp && baze);
	assign phi_out = bude;
	assign nphi    = dova;

	wire bele, atez, byju, alyp, buty, baly, afar, buvu, boga, asol, boma, byxo, bowa, afer, avor, alur;
	wire boga1mhz;
	dffr dffr_afer(boma, nt1_nt2, asol, afer); // check clk edge
	assign #T_INV  bele = !buto;
	assign #T_INV  atez = !clkin_a;
	assign #T_OR   byju = bele || atez;
	assign #T_INV  alyp = !taba;
	assign #T_INV  buty = !abol;
	assign #T_INV  baly = !byju;
	assign #T_NOR  afar = !(alyp || reset);
	assign #T_AND  buvu = buty && baly;
	assign #T_INV  boga = !baly;
	assign #T_OR   asol = afar || reset;
	assign #T_INV  byxo = !buvu;
	assign #T_INV  boma = !boga;
	assign #T_INV  bedo = !byxo;
	assign #T_INV  bowa = !bedo;
	assign #T_OR   avor = afer || asol;
	assign #T_INV  alur = !avor;
	assign boga1mhz = boga;
	assign to_cpu   = bowa;
	assign nreset2  = alur;

	wire tape, ufol, nreset_div;
	assign #T_AND  tape = ff04_ff07 && cpu_wr && tola_na1 && tovy_na0;
	assign #T_NOR  ufol = !(nclkin_a || reset || tape);
	assign nreset_div = ufol;

	wire tama, unyk, tero, uner, ufor, ukup, uvyn, tama16384;
	wire _16384hz, _32768hz, _65536hz, _131072hz, _262144hz, _524288hz;
	dffr dffr_tama(!unyk,    nreset_div, !tama, tama);
	dffr dffr_unyk(!tero,    nreset_div, !unyk, unyk);
	dffr dffr_tero(!uner,    nreset_div, !tero, tero);
	dffr dffr_uner(!ufor,    nreset_div, !uner, uner);
	dffr dffr_ufor(!ukup,    nreset_div, !ufor, ufor);
	dffr dffr_ukup(boga1mhz, nreset_div, !ukup, ukup);
	assign #T_INV  uvyn = !tama;
	assign tama16384 = !tama;
	assign _16384hz  = uvyn;
	assign _32768hz  = unyk;
	assign _65536hz  = tero;
	assign _131072hz = uner;
	assign _262144hz = ufor;
	assign _524288hz = ukup;

	wire ulur, ugot, tulu, tugo, tofe, teru, sola, subu, teka, uket, upof;
	wire umek, urek, utok, sapy, umer, rave, ryso, udor;
	wire tagy, tawu, taku, temu, tuse, upug, sepu, sawa, tatu;
	wire upyf, tubo, unut, taba, nff04_d0, nff04_d1;
	dffr dffr_ugot(ulur,  nreset_div, !ugot, ugot);
	dffr dffr_tulu(!ugot, nreset_div, !tulu, tulu);
	dffr dffr_tugo(!tulu, nreset_div, !tugo, tugo);
	dffr dffr_tofe(!tugo, nreset_div, !tofe, tofe);
	dffr dffr_teru(!tofe, nreset_div, !teru, teru);
	dffr dffr_sola(!teru, nreset_div, !sola, sola);
	dffr dffr_subu(!sola, nreset_div, !subu, subu);
	dffr dffr_teka(!subu, nreset_div, !teka, teka);
	dffr dffr_uket(!teka, nreset_div, !uket, uket);
	dffr dffr_upof(!uket, nreset_div, !upof, upof);
	assign #T_MUX  ulur = ff60_d1 ? boga1mhz : tama16384;
	assign #T_INV  umek = !ugot;
	assign #T_INV  urek = !tulu;
	assign #T_INV  utok = !tugo;
	assign #T_INV  sapy = !tofe;
	assign #T_INV  umer = !teru;
	assign #T_INV  rave = !sola;
	assign #T_INV  ryso = !subu;
	assign #T_INV  udor = !teka;
	assign #T_AND  tagy = ff04_ff07 && cpu_rd && tola_na1 && tovy_na0;
	assign #T_OR   upyf = reset || nclkin_a;
	assign #T_OR   tubo = clk_from_cpu || upyf;
	assign #T_AND  unut = upof && tubo;
	assign #T_OR   taba = nt1_t2 || t1_nt2 || unut;
	assign #T_TRI  tawu = tagy ? !umek : 1'bz;
	assign #T_TRI  taku = tagy ? !urek : 1'bz;
	assign #T_TRI  temu = tagy ? !utok : 1'bz;
	assign #T_TRI  tuse = tagy ? !sapy : 1'bz;
	assign #T_TRI  upug = tagy ? !umer : 1'bz;
	assign #T_TRI  sepu = tagy ? !rave : 1'bz;
	assign #T_TRI  sawa = tagy ? !ryso : 1'bz;
	assign #T_TRI  tatu = tagy ? !udor : 1'bz;
	assign nff04_d0 = umek;
	assign nff04_d1 = urek;
	assign d = { tatu, sawa, sepu, upug, tuse, temu, taku, tawu };

	wire atus, coke, bara, caru, bylu, bure, fyne, culo, apef, gale, beze, bule, gexy, cofu, baru, horu, bufy, byfe;
	wire _512hz, _256hz, _128hz, horu_512hz, bufy_256hz;
	dffr dffr_bara(coke,  atus, umer,  bara); // check edge
	dffr dffr_caru(bure,  atus, !caru, caru); // check edge
	dffr dffr_bylu(!caru, atus, !bylu, bylu); // check edge
	assign #T_INV  atus = !apu_reset;
	assign #T_INV  coke = !ajer_2mhz;
	assign #T_INV  bure = bara; /* takes !q output of dff */
	assign #T_INV  fyne = !bure;
	assign #T_INV  culo = caru; /* takes !q output of dff */
	assign #T_INV  apef = bylu; /* takes !q output of dff */
	assign #T_MUX  gale = fero_q ? hama_512k : fyne;
	assign #T_MUX  beze = fero_q ? hama_512k : culo;
	assign #T_MUX  bule = fero_q ? hama_512k : apef;
	assign #T_INV  gexy = !gale;
	assign #T_INV  horu = !gexy;
	assign #T_INV  cofu = !beze;
	assign #T_INV  bufy = !cofu;
	assign #T_INV  baru = !bule;
	assign #T_INV  byfe = !baru;
	assign _512hz = bara;
	assign _256hz = caru;
	assign _128hz = bylu;
	assign horu_512hz = horu;
	assign bufy_256hz = bufy;
	assign byfe_128hz = byfe;

	wire bopo, atyk, avok, bavu, jeso, hama, bavu_1mhz, _2097152hz, _1048576hz, jeso_512k, hama_512k;
	dffr dffr_atyk(aryf_4mhz, bopo,        !atyk, atyk); // check edge
	dffr dffr_avok(atyk,      bopo,        !avok, avok); // check edge
	dffr dffr_jeso(bavu,      napu_reset5, !jeso, jeso); // check edge
	assign #T_INV  bopo = !apu_reset;
	assign #T_INV  bavu = !avok;
	assign #T_INV  hama = jeso; /* takes !q output of dff */
	assign _2097152hz = atyk;
	assign _1048576hz = avok;
	assign jeso_512k = jeso;
	assign hama_512k = hama;

endmodule

module dma(
		clk1, d, ma, dma_a,
		nreset6, from_cpu5,
		cpu_rd2, cpu_wr2, ff46,
		amab, wyja, caty, dma_run,
		vram_to_oam, dma_addr_ext, oam_addr_dma,
		nphi_out, mopa_phi
	);

	inout  wire [7:0] d;
	output wire [12:0] ma;
	output wire [15:0] dma_a;

	input wire clk1, nreset6, from_cpu5;
	input wire cpu_rd2, cpu_wr2, ff46;

	input  wire amab, nphi_out;
	output wire wyja, caty, dma_run, mopa_phi;
	output wire vram_to_oam, dma_addr_ext, oam_addr_dma;

	wire decy, maka, naxy, powu, luvy, molu, nygo, pusy, lavy, loru, lyxe, lupa, ahoc, loko, lapa, meta;
	dffr dffr_maka(clk1,     nreset6, caty, maka); // check edge
	dffr dffr_luvy(nphi_out, nreset6, lupa, luvy); // check edge
	assign #T_INV  decy = !from_cpu5;
	assign #T_INV  caty = !decy;
	assign #T_NOR  naxy = !(maka || luvy);
	assign #T_AND  powu = matu && naxy;
	assign #T_AO   wyja = (amab && cpu_wr2) || powu;
	assign #T_AND  molu = ff46 && cpu_rd2;
	assign #T_INV  nygo = !molu;
	assign #T_INV  pusy = !nygo;
	assign #T_AND  lavy = ff46 && cpu_wr2;
	assign #T_INV  loru = !lavy;
	assign #T_OR   lyxe = loru || loko;
	assign #T_NOR  lupa = !(lavy || lyxe);
	assign #T_INV  ahoc = !vram_to_oam;
	assign #T_NAND loko = !(nreset6 && !lene);
	assign #T_INV  lapa = !loko;
	assign #T_AND  meta = nphi_out && loky;

	wire mopa, navo, nolo, myte, lene, lara, loky, matu, mory, luma, logo, duga, lebu, muda, muho, lufa;
	dffr dffr_myte(mopa,     lapa,    nolo, myte); // check edge
	dffr dffr_lene(mopa,     nreset6, luvy, lene); // check edge
	dffr dffr_matu(nphi_out, nreset6, loky, matu); // check edge
	assign #T_INV  mopa = !nphi_out;
	assign #T_NAND navo = !(dma_a[0] && dma_a[1] && dma_a[2] && dma_a[3] && dma_a[4] && dma_a[7]);
	assign #T_INV  nolo = !navo;
	assign #T_NAND lara = !(loky && !myte && nreset6);
	assign #T_NAND loky = !(lara && !lene);
	assign #T_NAND mory = !(matu && logo);
	assign #T_INV  luma = !mory;
	assign #T_INV  logo = !muda;
	assign #T_INV  duga = !matu;
	assign #T_INV  lebu = !dma_a[15];
	assign #T_NOR  muda = !(dma_a[13] || dma_a[14] || lebu);
	assign #T_NAND muho = !(matu && muda);
	assign #T_INV  lufa = !muho;
	assign mopa_phi     = mopa;
	assign dma_run      = matu;
	assign dma_addr_ext = luma;
	assign oam_addr_dma = duga;
	assign vram_to_oam  = lufa;

	wire nafa, nygy, para, pyne, pula, nydo, poku, maru, poly, pare, rema, rofo, raly, pane, resu, nuvy;
	wire evax, exyf, eraf, duve, fusy;
	dff dff_nafa(loru, d[0], nafa); // check edge
	dff dff_nygy(loru, d[4], nygy); // check edge
	dff dff_para(loru, d[2], para); // check edge
	dff dff_pyne(loru, d[1], pyne); // check edge
	dff dff_pula(loru, d[5], pula); // check edge
	dff dff_nydo(loru, d[3], nydo); // check edge
	dff dff_poku(loru, d[6], poku); // check edge
	dff dff_maru(loru, d[7], maru); // check edge
	assign #T_TRI  poly = pusy ? nafa : 1'bz; /* takes !q output of dff */
	assign #T_TRI  pare = pusy ? nygy : 1'bz; /* takes !q output of dff */
	assign #T_TRI  rema = pusy ? para : 1'bz; /* takes !q output of dff */
	assign #T_TRI  rofo = pusy ? pyne : 1'bz; /* takes !q output of dff */
	assign #T_TRI  raly = pusy ? pula : 1'bz; /* takes !q output of dff */
	assign #T_TRI  pane = pusy ? nydo : 1'bz; /* takes !q output of dff */
	assign #T_TRI  resu = pusy ? poku : 1'bz; /* takes !q output of dff */
	assign #T_TRI  nuvy = pusy ? maru : 1'bz; /* takes !q output of dff */
	assign #T_TRI  evax = !ahoc ? !nafa : 1'bz;
	assign #T_TRI  exyf = !ahoc ? !nygy : 1'bz;
	assign #T_TRI  eraf = !ahoc ? !para : 1'bz;
	assign #T_TRI  duve = !ahoc ? !pyne : 1'bz;
	assign #T_TRI  fusy = !ahoc ? !nydo : 1'bz;
	assign d[0] = poly;
	assign d[4] = pare;
	assign d[2] = rema;
	assign d[1] = rofo;
	assign d[5] = raly;
	assign d[3] = pane;
	assign d[6] = resu;
	assign d[7] = nuvy;
	assign dma_a[8]  = nafa;
	assign dma_a[12] = nygy;
	assign dma_a[10] = para;
	assign dma_a[9]  = pyne;
	assign dma_a[13] = pula;
	assign dma_a[11] = nydo;
	assign dma_a[14] = poku;
	assign dma_a[15] = maru;
	assign ma[8]  = evax;
	assign ma[12] = exyf;
	assign ma[10] = eraf;
	assign ma[9]  = duve;
	assign ma[11] = fusy;

	wire naky, pyro, nefy, muty, nyko, pylo, nuto, mugu, ecal, egez, fuhe, fyzy, damu, dava, eteg, erew;
	dffr dffr_naky(meta,  lapa, !naky, naky); // check edge
	dffr dffr_pyro(!naky, lapa, !pyro, pyro); // check edge
	dffr dffr_nefy(!pyro, lapa, !nefy, nefy); // check edge
	dffr dffr_muty(!nefy, lapa, !muty, muty); // check edge
	dffr dffr_nyko(!muty, lapa, !nyko, nyko); // check edge
	dffr dffr_pylo(!nyko, lapa, !pylo, pylo); // check edge
	dffr dffr_nuto(!pylo, lapa, !nuto, nuto); // check edge
	dffr dffr_mugu(!nuto, lapa, !mugu, mugu); // check edge
	assign #T_TRI  ecal = !ahoc ? !naky : 1'bz;
	assign #T_TRI  egez = !ahoc ? !pyro : 1'bz;
	assign #T_TRI  fuhe = !ahoc ? !nefy : 1'bz;
	assign #T_TRI  fyzy = !ahoc ? !muty : 1'bz;
	assign #T_TRI  damu = !ahoc ? !nyko : 1'bz;
	assign #T_TRI  dava = !ahoc ? !pylo : 1'bz;
	assign #T_TRI  eteg = !ahoc ? !nuto : 1'bz;
	assign #T_TRI  erew = !ahoc ? !mugu : 1'bz;
	assign dma_a[0] = naky;
	assign dma_a[1] = pyro;
	assign dma_a[2] = nefy;
	assign dma_a[3] = muty;
	assign dma_a[4] = nyko;
	assign dma_a[5] = pylo;
	assign dma_a[6] = nuto;
	assign dma_a[7] = mugu;
	assign ma[0] = ecal;
	assign ma[1] = egez;
	assign ma[2] = fuhe;
	assign ma[3] = fyzy;
	assign ma[4] = damu;
	assign ma[5] = dava;
	assign ma[6] = eteg;
	assign ma[7] = erew;

endmodule

module sys_decode(
		reset, nreset2, t1, t2, wr_in, rd_b, a, d,
		cpu_rd_sync, cpu_raw_rd, cpu_wr_raw,
		from_cpu6, to_cpu_tutu,
		cpu_wr, cpu_wr2, cpu_rd, cpu_rd2,
		nt1_nt2, nt1_t2, t1_nt2,
		ff04_ff07, ff0f_rd, ff0f_wr,
		hram_cs,
		anap, bedo, tutu,
		a00_07, ffxx, nffxx, nfexxffxx, saro,
		ff60_d1, ff60_d0, boot_cs
	);

	input  wire reset, nreset2, t1, t2, wr_in, rd_b;
	input  wire [15:0] a;
	inout  wire [7:0] d;
	input  wire cpu_rd_sync, cpu_raw_rd, cpu_wr_raw;
	input  wire from_cpu6;
	output wire to_cpu_tutu;
	output wire cpu_wr, cpu_wr2, cpu_rd, cpu_rd2;
	output wire nt1_nt2, nt1_t2, t1_nt2;

	output wire ff04_ff07, ff0f_rd, ff0f_wr;
	output wire hram_cs;

	input  wire anap, bedo;
	output wire tutu;
	input  wire a00_07;
	output wire ffxx, nffxx, nfexxffxx, saro;
	output wire ff60_d1, ff60_d0;
	output wire boot_cs;

	wire ubet, uvar, upoj, unor, umut;
	assign #T_INV  ubet = !t1;
	assign #T_INV  uvar = !t2;
	assign #T_NAND upoj = !(ubet && uvar && reset);
	assign #T_AND  unor = t2 && ubet;
	assign #T_AND  umut = uvar && t1;
	assign nt1_nt2 = upoj;
	assign nt1_t2  = unor;
	assign t1_nt2  = umut;

	wire ubal, ujyv, lexy, tapu, tedo, dyky, ajas, cupa, asot, pin_nc;
	assign #T_MUX  ubal = !(nt1_t2 ? wr_in : cpu_rd_sync);
	assign #T_MUX  ujyv = !(nt1_t2 ? rd_b  : cpu_raw_rd);
	assign #T_INV  lexy = !from_cpu6;
	assign #T_INV  tapu = !ubal;
	assign #T_INV  tedo = !ujyv;
	assign #T_INV  dyky = !tapu;
	assign #T_INV  ajas = !tedo;
	assign #T_INV  cupa = !dyky;
	assign #T_INV  asot = !ajas;
	assign pin_nc  = lexy;
	assign cpu_wr  = tapu;
	assign cpu_wr2 = cupa;
	assign cpu_rd  = tedo;
	assign cpu_rd2 = asot;

	wire ryfo, semy, sapa, rolo, refa;
	assign #T_AND  ryfo = a[2] && a00_07 && ffxx;
	assign #T_NOR  semy = !(a[7] || a[6] || a[5] || a[4]);
	assign #T_AND  sapa = a[0] && a[1] && a[2] && a[3];
	assign #T_NAND rolo = !(semy && sapa && ffxx && cpu_rd);
	assign #T_NAND refa = !(semy && sapa && ffxx && cpu_wr_raw);
	assign ff04_ff07 = ryfo;
	assign ff0f_rd   = rolo;
	assign ff0f_wr   = refa;

	wire zyra, zage, zabu, zoke, zera, zufy, zyky, zyga, zovy, zuko, zuvy, zyba, zole, zaje, zubu, zapy;
	wire zete, zefu, zyro, zapa, bootrom_na7, bootrom_na6, bootrom_na3, bootrom_na2;
	wire bootrom_na5_na4, bootrom_na5_a4, bootrom_a5_na4, bootrom_a5_a4;
	wire bootrom_na1_na0, bootrom_na1_a0, bootrom_a1_na0, bootrom_a1_a0;
	assign #T_INV  zyra = !a[7];
	assign #T_INV  zage = !a[6];
	assign #T_INV  zabu = !a[3];
	assign #T_INV  zoke = !a[2];
	assign #T_INV  zera = !a[5];
	assign #T_INV  zufy = !a[4];
	assign #T_AND  zyky = zera && zufy;
	assign #T_AND  zyga = zera && a[4];
	assign #T_AND  zovy = a[5] && zufy;
	assign #T_AND  zuko = a[5] && a[4];
	assign #T_INV  zuvy = !a[1];
	assign #T_INV  zyba = !a[0];
	assign #T_AND  zole = zuvy && zyba;
	assign #T_AND  zaje = zuvy && a[0];
	assign #T_AND  zubu = zyba && a[1];
	assign #T_AND  zapy = a[1] && a[0];
	assign #T_INV  zete = !zole;
	assign #T_INV  zefu = !zaje;
	assign #T_INV  zyro = !zubu;
	assign #T_INV  zapa = !zapy;
	assign bootrom_na7     = zyra;
	assign bootrom_na6     = zage;
	assign bootrom_na3     = zabu;
	assign bootrom_na2     = zoke;
	assign bootrom_na5_na4 = zyky;
	assign bootrom_na5_a4  = zyga;
	assign bootrom_a5_na4  = zovy;
	assign bootrom_a5_a4   = zuko;
	assign bootrom_na1_na0 = zete;
	assign bootrom_na1_a0  = zefu;
	assign bootrom_a1_na0  = zyro;
	assign bootrom_a1_a0   = zapa;

	wire apet, aper, amut, buro;
	assign #T_OR   apet = nt1_t2 || t1_nt2;
	assign #T_NAND aper = !(apet && a[5] && a[6] && cpu_wr && anap);
	dffr dffr_amut(aper, nreset2, d[1], amut); // check edge
	dffr dffr_buro(aper, nreset2, d[0], buro); // check edge
	assign ff60_d1 = amut;
	assign ff60_d0 = buro;

	wire leco, raru, rowe, ryke, ryne, rase, rejy, reka, romy;
	assign #T_NOR  leco = !(bedo || nt1_t2);
	assign #T_TRI  raru = leco ? 1'b1 : 1'bz;
	assign #T_TRI  rowe = leco ? 1'b1 : 1'bz;
	assign #T_TRI  ryke = leco ? 1'b1 : 1'bz;
	assign #T_TRI  ryne = leco ? 1'b1 : 1'bz;
	assign #T_TRI  rase = leco ? 1'b1 : 1'bz;
	assign #T_TRI  rejy = leco ? 1'b1 : 1'bz;
	assign #T_TRI  reka = leco ? 1'b1 : 1'bz;
	assign #T_TRI  romy = leco ? 1'b1 : 1'bz;
	assign d[7] = raru;
	assign d[5] = rowe;
	assign d[6] = ryke;
	assign d[1] = ryne;
	assign d[3] = rase;
	assign d[2] = rejy;
	assign d[4] = reka;
	assign d[0] = romy;

	wire wale, woly, wuta;
	assign #T_NAND wale = !(a[0] && a[1] && a[2] && a[3] && a[4] && a[5] && a[6]);
	assign #T_NAND woly = !(wale && a[7] && ffxx);
	assign #T_INV  wuta = !woly;
	assign hram_cs = woly;

	wire tona, syke, bako, tuna, rycu, rope, soha;
	assign #T_INV  tona = !a[8];
	assign #T_NAND tuna = !(a[15] && a[14] && a[13] && a[12] && a[11] && a[10] && a[9]);
	assign #T_NOR  syke = !(tona || tuna);
	assign #T_INV  bako = !syke;
	assign #T_INV  rycu = !tuna;
	assign #T_INV  soha = !ffxx;
	assign #T_NAND rope = !(rycu && soha);
	assign #T_INV  saro = !rope;
	assign ffxx      = syke;
	assign nffxx     = bako;
	assign nfexxffxx = tuna;

	wire tyro, tufa, texe, sato, tuge, tepu, sypu, tera, yaza, yula, tulo, zoro, zadu, zufa, zado, zery;
	dffr dffr_tepu(tuge, nreset2, sato, tepu); // check edge
	assign #T_NOR  tyro = !(a[7] || a[5] || a[3] || a[2] || a[1] || a[0]);
	assign #T_AND  tufa = a[4] && a[6];
	assign #T_AND  texe = cpu_rd && ffxx && tufa && tyro;
	assign #T_OR   sato = d[0] || tepu;
	assign #T_NAND tuge = !(tyro && tufa && ffxx && cpu_wr);
	assign #T_TRI  sypu = texe ? tepu : 1'bz; /* takes !q output of dff */
	assign #T_INV  tera = !tepu;
	assign #T_INV  yaza = t1_nt2;
	assign #T_AND  tutu = tera && tulo;
	assign #T_AND  yula = yaza && tutu && cpu_rd;
	assign #T_NOR  tulo = !(a[15] || a[14] || a[13] || a[12] || a[11] || a[10] || a[9] || a[8]);
	assign #T_NOR  zoro = !(a[15] || a[14] || a[13] || a[12]);
	assign #T_NOR  zadu = !(a[11] || a[10] || a[9] || a[8]);
	assign #T_AND  zufa = zoro && zadu;
	assign #T_NAND zado = !(yula && zufa);
	assign #T_INV  zery = !zado;
	assign to_cpu_tutu = tutu;
	assign boot_cs     = zery;

endmodule

module ext_cpu_busses(
		d, d_in, d_d,
		a, a_c, a_a, a_d, dma_a,
		wr_a, wr_c, rd_a, rd_c,
		from_cpu3, from_cpu4, from_cpu5,
		cpu_raw_rd, cpu_rd_sync,
		cpu_rd, t1_nt2, nt1_t2, dma_addr_ext,
		abuz, tutu, texo, roru, lula, nfexxffxx,
		ncs_out, tola_na1
	);

	inout  wire [7:0]  d;
	input  wire [7:0]  d_in;
	output wire [7:0]  d_d;
	inout  wire [15:0] a;
	input  wire [15:0] a_c, dma_a;
	output wire [15:0] a_a, a_d;

	output wire wr_a, wr_c, rd_a, rd_c;

	input wire from_cpu3, from_cpu4, from_cpu5;
	input wire cpu_raw_rd, cpu_rd_sync;
	input wire cpu_rd, t1_nt2, nt1_t2, dma_addr_ext;

	input  wire abuz, tutu, nfexxffxx;
	output wire texo, roru, lula;

	output wire ncs_out, tola_na1;

	wire sogy, tuma, tynu, toza, soby, sepy, ryca, raza, syzu, tyho, tazy, rulo, suze;
	assign #T_INV  sogy = !a[14];
	assign #T_AND  tuma = a[13] && sogy && a[15];
	assign #T_AO   tynu = (a[15] && a[14]) || tuma;
	assign #T_AND  toza = tynu && abuz && nfexxffxx;
	assign #T_NOR  soby = !(a[15] || tutu);
	assign #T_NAND sepy = !(abuz && soby);
	assign #T_INV  ryca = !nt1_t2;
	assign #T_INV  raza = a_c[15];
	assign #T_TRI  syzu = !ryca ? !raza : 1'bz;
	assign #T_MUX  tyho = dma_addr_ext ? dma_a[15] : toza;
	assign #T_MUX  tazy = dma_addr_ext ? dma_a[15] : sepy;
	assign #T_NOR  rulo = !(nt1_t2 || tazy);
	assign #T_NAND suze = !(tazy && ryca);
	assign ncs_out = tyho;
	assign a_d[15] = rulo;
	assign a_a[15] = suze;
	assign a[15]   = syzu;

	wire tova, nyre, lonu, lobu, lumy, pate, lysa, luno, pege, muce, mojy, male, pamy, masu, mano;
	wire pahy, puhe, leva, labe, loso, luce, lyny, lepy, rore, roxu, meny, mune, mego, myny, net01;
	latch latch_nyre(mate, a[14], nyre);
	latch latch_lonu(mate, a[13], lonu);
	latch latch_lobu(mate, a[12], lobu);
	latch latch_lumy(mate, a[11], lumy);
	latch latch_pate(mate, a[10], pate);
	latch latch_lysa(mate, a[9],  lysa);
	latch latch_luno(mate, a[8],  luno);
	assign #T_INV  tova = !nt1_t2;
	assign #T_MUX  pege = dma_addr_ext ? dma_a[14] : nyre;
	assign #T_MUX  muce = dma_addr_ext ? dma_a[13] : lonu;
	assign #T_MUX  mojy = dma_addr_ext ? dma_a[12] : lobu;
	assign #T_MUX  male = dma_addr_ext ? dma_a[11] : lumy;
	assign #T_MUX  pamy = dma_addr_ext ? dma_a[10] : pate;
	assign #T_MUX  masu = dma_addr_ext ? dma_a[9]  : lysa;
	assign #T_MUX  mano = dma_addr_ext ? dma_a[8]  : luno;
	assign #T_NOR  pahy = !(nt1_t2 || pege);
	assign #T_NAND puhe = !(pege && tova);
	assign #T_NOR  leva = !(nt1_t2 || muce);
	assign #T_NAND labe = !(muce && tova);
	assign #T_NOR  loso = !(nt1_t2 || mojy);
	assign #T_NAND luce = !(mojy && tova);
	assign #T_NOR  lyny = !(nt1_t2 || male);
	assign #T_NAND lepy = !(male && tova);
	assign #T_NOR  rore = !(nt1_t2 || pamy);
	assign #T_NAND roxu = !(pamy && tova);
	assign #T_NOR  meny = !(nt1_t2 || masu);
	assign #T_NAND mune = !(masu && tova);
	assign #T_NOR  mego = !(nt1_t2 || mano);
	assign #T_NAND myny = !(mano && tova);
	assign net01   = tova;
	assign a_d[14] = pahy;
	assign a_a[14] = puhe;
	assign a_d[13] = leva;
	assign a_a[13] = labe;
	assign a_d[12] = loso;
	assign a_a[12] = luce;
	assign a_d[11] = lyny;
	assign a_a[11] = lepy;
	assign a_d[10] = rore;
	assign a_a[10] = roxu;
	assign a_d[9]  = meny;
	assign a_a[9]  = mune;
	assign a_d[8]  = mego;
	assign a_a[8]  = myny;

	wire arym, aros, atev, avys, aret, alyr, apur, alor, asur, atyr, atov, atem, amer, apok, atol, amet;
	wire colo, defy, cyka, cepu, ajav, badu, bevo, byla, bola, boty, bajo, boku, cotu, caba, koty, kupo;
	latch latch_arym(mate, a[7], arym);
	latch latch_aros(mate, a[6], aros);
	latch latch_atev(mate, a[5], atev);
	latch latch_avys(mate, a[4], avys);
	latch latch_aret(mate, a[3], aret);
	latch latch_alyr(mate, a[2], alyr);
	latch latch_apur(mate, a[1], apur);
	latch latch_alor(mate, a[0], alor);
	assign #T_MUX  asur = dma_addr_ext ? dma_a[7] : arym;
	assign #T_MUX  atyr = dma_addr_ext ? dma_a[6] : aros;
	assign #T_MUX  atov = dma_addr_ext ? dma_a[5] : atev;
	assign #T_MUX  atem = dma_addr_ext ? dma_a[4] : avys;
	assign #T_MUX  amer = dma_addr_ext ? dma_a[3] : aret;
	assign #T_MUX  apok = dma_addr_ext ? dma_a[2] : alyr;
	assign #T_MUX  atol = dma_addr_ext ? dma_a[1] : apur;
	assign #T_MUX  amet = dma_addr_ext ? dma_a[0] : alor;
	assign #T_NOR  colo = !(nt1_t2 || asur);
	assign #T_NAND defy = !(net01 && asur);
	assign #T_NOR  cyka = !(nt1_t2 || atyr);
	assign #T_NAND cepu = !(net01 && atyr);
	assign #T_NOR  ajav = !(nt1_t2 || atov);
	assign #T_NAND badu = !(net01 && atov);
	assign #T_NOR  bevo = !(nt1_t2 || atem);
	assign #T_NAND byla = !(net01 && atem);
	assign #T_NOR  bola = !(nt1_t2 || amer);
	assign #T_NAND boty = !(net01 && amer);
	assign #T_NOR  bajo = !(nt1_t2 || apok);
	assign #T_NAND boku = !(net01 && apok);
	assign #T_NOR  cotu = !(nt1_t2 || atol);
	assign #T_NAND caba = !(net01 && atol);
	assign #T_NOR  koty = !(nt1_t2 || amet);
	assign #T_NAND kupo = !(net01 && amet);
	assign a_d[7] = colo;
	assign a_a[7] = defy;
	assign a_d[6] = cyka;
	assign a_a[6] = cepu;
	assign a_d[5] = ajav;
	assign a_a[5] = badu;
	assign a_d[4] = bevo;
	assign a_a[4] = byla;
	assign a_d[3] = bola;
	assign a_a[3] = boty;
	assign a_d[2] = bajo;
	assign a_a[2] = boku;
	assign a_d[1] = cotu;
	assign a_a[1] = caba;
	assign a_d[0] = koty;
	assign a_a[0] = kupo;

	wire tola, mule, loxo, lasy, mate, sore, tevy, levo, lagu;
	assign #T_INV  tola = !a[1];
	assign #T_INV  mule = !t1_nt2;
	assign #T_AO   loxo = (mule && texo) || t1_nt2;
	assign #T_INV  lasy = !loxo;
	assign #T_INV  mate = !lasy;
	assign #T_INV  sore = !a[15];
	assign #T_OR   tevy = a[13] || a[14] || sore;
	assign #T_AND  texo = from_cpu4 && tevy;
	assign #T_INV  levo = !texo;
	assign #T_AO   lagu = (cpu_raw_rd && levo) || from_cpu3;
	assign tola_na1 = tola;

	wire moca, mexo, lywe, nevy, moty, puva, tymu, usuf, uver, ugac, urun;
	assign #T_NOR  moca = !(texo || t1_nt2);
	assign #T_INV  mexo = !cpu_rd_sync;
	assign #T_INV  lywe = !lagu;
	assign #T_OR   nevy = mexo || moca;
	assign #T_OR   moty = moca || lywe;
	assign #T_OR   puva = nevy || dma_addr_ext;
	assign #T_NOR  tymu = !(dma_addr_ext || moty);
	assign #T_NOR  usuf = !(nt1_t2 || puva);
	assign #T_NAND uver = !(puva && net01);
	assign #T_NAND ugac = !(net01 && tymu);
	assign #T_NOR  urun = !(tymu || nt1_t2);
	assign wr_c = usuf;
	assign wr_a = uver;
	assign rd_a = ugac;
	assign rd_c = urun;

	wire base, afec, buxu, camu, cygu, cogo, kova, anar, azuv, akan, byxe, byne, byna, kejo;
	assign #T_INV  base = !a_c[3];
	assign #T_INV  afec = !a_c[4];
	assign #T_INV  buxu = !a_c[2];
	assign #T_INV  camu = !a_c[1];
	assign #T_INV  cygu = !a_c[6];
	assign #T_INV  cogo = !a_c[7];
	assign #T_INV  kova = !a_c[0];
	assign #T_TRI  anar = !net01 ? !base : 1'bz;
	assign #T_TRI  azuv = !net01 ? !afec : 1'bz;
	assign #T_TRI  akan = !net01 ? !buxu : 1'bz;
	assign #T_TRI  byxe = !net01 ? !camu : 1'bz;
	assign #T_TRI  byne = !net01 ? !cygu : 1'bz;
	assign #T_TRI  byna = !net01 ? !cogo : 1'bz;
	assign #T_TRI  kejo = !net01 ? !kova : 1'bz;
	assign a[3] = anar;
	assign a[4] = azuv;
	assign a[2] = akan;
	assign a[1] = byxe;
	assign a[6] = byne;
	assign a[7] = byna;
	assign a[0] = kejo;

	wire lahe, lura, mujy, pevo, mady, nena, sura, abup, lyna, lefy, lofa, nefe, lora, mapu, rala, ajov;
	assign #T_INV  lahe = !a_c[12];
	assign #T_INV  lura = !a_c[13];
	assign #T_INV  mujy = !a_c[8];
	assign #T_INV  pevo = !a_c[14];
	assign #T_INV  mady = !a_c[11];
	assign #T_INV  nena = !a_c[9];
	assign #T_INV  sura = !a_c[10];
	assign #T_INV  abup = !a_c[5];
	assign #T_TRI  lyna = !net01 ? !lahe : 1'bz;
	assign #T_TRI  lefy = !net01 ? !lura : 1'bz;
	assign #T_TRI  lofa = !net01 ? !mujy : 1'bz;
	assign #T_TRI  nefe = !net01 ? !pevo : 1'bz;
	assign #T_TRI  lora = !net01 ? !mady : 1'bz;
	assign #T_TRI  mapu = !net01 ? !nena : 1'bz;
	assign #T_TRI  rala = !net01 ? !sura : 1'bz;
	assign #T_TRI  ajov = !net01 ? !abup : 1'bz;
	assign a[12] = lyna;
	assign a[13] = lefy;
	assign a[8]  = lofa;
	assign a[14] = nefe;
	assign a[11] = lora;
	assign a[9]  = mapu;
	assign a[10] = rala;
	assign a[5]  = ajov;

	wire redu, rogy, ryda, rune, resy, rypu, suly, seze, tamu;
	assign #T_INV  redu = !cpu_rd;
	assign #T_MUX  roru = nt1_t2 ? redu : moty;
	assign #T_INV  lula = !roru;
	assign #T_NOR  rogy = !(roru || d[6]);
	assign #T_NOR  ryda = !(roru || d[7]);
	assign #T_NOR  rune = !(roru || d[0]);
	assign #T_NOR  resy = !(roru || d[4]);
	assign #T_NOR  rypu = !(roru || d[1]);
	assign #T_NOR  suly = !(roru || d[2]);
	assign #T_NOR  seze = !(roru || d[3]);
	assign #T_NOR  tamu = !(roru || d[5]);
	assign d_d[6] = rogy;
	assign d_d[7] = ryda;
	assign d_d[0] = rune;
	assign d_d[4] = resy;
	assign d_d[1] = rypu;
	assign d_d[2] = suly;
	assign d_d[3] = seze;
	assign d_d[5] = tamu;

	wire lavo, sody, selo, rony, soma, raxy, rupa, sago, sazy;
	wire tepe, tavo, ruvo, ryma, ryko, sevu, safo, taju;
	latch latch_sody(lavo, d_in[4], sody);
	latch latch_selo(lavo, d_in[3], selo);
	latch latch_rony(lavo, d_in[1], rony);
	latch latch_soma(lavo, d_in[0], soma);
	latch latch_raxy(lavo, d_in[2], raxy);
	latch latch_rupa(lavo, d_in[6], rupa);
	latch latch_sago(lavo, d_in[5], sago);
	latch latch_sazy(lavo, d_in[7], sazy);
	assign #T_NAND lavo = !(cpu_raw_rd && texo && from_cpu5);
	assign #T_TRI  tepe = !lavo ? !sody : 1'bz;
	assign #T_TRI  tavo = !lavo ? !selo : 1'bz;
	assign #T_TRI  ruvo = !lavo ? !rony : 1'bz;
	assign #T_TRI  ryma = !lavo ? !soma : 1'bz;
	assign #T_TRI  ryko = !lavo ? !raxy : 1'bz;
	assign #T_TRI  sevu = !lavo ? !rupa : 1'bz;
	assign #T_TRI  safo = !lavo ? !sago : 1'bz;
	assign #T_TRI  taju = !lavo ? !sazy : 1'bz;
	assign d[4] = tepe;
	assign d[3] = tavo;
	assign d[1] = ruvo;
	assign d[0] = ryma;
	assign d[2] = ryko;
	assign d[6] = sevu;
	assign d[5] = safo;
	assign d[7] = taju;

endmodule

module apu_ctrl(
		cpu_rd, ncpu_rd,
		nreset2,
		d,
		from_cpu,
		ff24, ff25, ff26,
		apu_wr,
		apu_reset, net03,
		napu_reset, napu_reset2, napu_reset4, napu_reset5, napu_reset6,
		apuv_4mhz, ajer_2mhz, byfe_128hz, dyfa_1mhz,
		fero_q, cate, gaxo,
		lmixer, rmixer,
		nch1_active, nch2_active, nch3_active, nch4_active
	);

	input wire cpu_rd;
	input wire nreset2;

	inout wire [7:0] d;

	input wire from_cpu;

	input wire ff24, ff25, ff26;

	input  wire apu_wr;
	output wire apu_reset, net03, ncpu_rd;
	output wire napu_reset, napu_reset2, napu_reset4, napu_reset5, napu_reset6;
	input  wire apuv_4mhz;
	output wire ajer_2mhz, dyfa_1mhz;
	input  wire byfe_128hz;
	output wire fero_q, cate, gaxo;

	output wire [3:0] lmixer, rmixer;

	input wire nch1_active, nch2_active, nch3_active, nch4_active;

	wire ajer, bata, calo, dyfa, najer_2mhz;
	dffr dffr_ajer(apuv_4mhz, napu_reset3, !ajer, ajer); // check edge
	dffr dffr_calo(bata,      napu_reset,  !calo, calo); // check edge
	assign #T_INV  bata = !ajer_2mhz;
	assign #T_INV  dyfa = calo; /* takes !q output of dff */
	assign ajer_2mhz  = ajer;
	assign najer_2mhz = !ajer;
	assign dyfa_1mhz  = dyfa;

	wire dapa, afat, agur, atyv, kame, cepo, napu_reset3;
	assign #T_INV  dapa = !apu_reset;
	assign #T_INV  afat = !apu_reset;
	assign #T_INV  agur = !apu_reset;
	assign #T_INV  atyv = !apu_reset;
	assign #T_INV  kame = !apu_reset;
	assign #T_INV  cepo = !apu_reset;
	assign napu_reset4 = dapa;
	assign napu_reset2 = afat;
	assign napu_reset  = agur;
	assign napu_reset3 = atyv;
	assign napu_reset5 = kame;
	assign napu_reset6 = cepo;

	wire kydu, jure, hapo, gufo, jyro, kuby, keba, hawu, hada, hope, bopy, bowy, baza, cely, cone;
	wire kepy, etuc, foku, efop, fero, edek;
	dffr dffr_hada(hawu,       gufo,        d[7], hada); // check edge
	dffr dffr_bowy(bopy,       kepy,        d[5], bowy); // check edge
	dffr dffr_baza(najer_2mhz, napu_reset3, bowy, baza); // check edge
	dffr dffr_fero(foku,       kepy,        efop, fero); // check edge
	assign #T_INV  kydu = !ncpu_rd;
	assign #T_NAND jure = !(kydu && ff26);
	assign #T_NAND hawu = !(ff26 && apu_wr);
	assign #T_NAND bopy = !(apu_wr && ff26);
	assign #T_INV  kepy = !jyro;
	assign #T_INV  hapo = !nreset2;
	assign #T_INV  gufo = !hapo;
	assign #T_OR   jyro = hapo || !hada;
	assign #T_TRI  hope = !jure ? !hada : 1'bz;
	assign #T_INV  kuby = !jyro;
	assign #T_INV  keba = !kuby;
	assign #T_MUX  cely = net03 ? baza : byfe_128hz;
	assign #T_INV  cone = !cely;
	assign #T_INV  cate = !cone;
	assign #T_AND  etuc = apu_wr && ff26;
	assign #T_AND  efop = d[4] && from_cpu;
	assign #T_INV  foku = !etuc;
	assign #T_INV  edek = fero; /* takes !q output of dff */
	assign apu_reset = keba;
	assign fero_q    = fero;
	assign net03     = edek;
	assign d[7]      = hope;

	wire aguz, byma, befu, adak, bosu, baxy, bubu, bowe, ataf;
	wire bedu, cozu, bumo, byre, apos, ager, byga, apeg;
	wire atum, bocy, arux, amad, axem, avud, awed, akod;
	dffr dffr_bedu(bubu, jyro, d[7], bedu); // check edge
	dffr dffr_cozu(bubu, jyro, d[6], cozu); // check edge
	dffr dffr_bumo(bubu, jyro, d[5], bumo); // check edge
	dffr dffr_byre(bubu, jyro, d[4], byre); // check edge
	dffr dffr_apos(ataf, jyro, d[3], apos); // check edge
	dffr dffr_ager(ataf, jyro, d[2], ager); // check edge
	dffr dffr_byga(ataf, jyro, d[1], byga); // check edge
	dffr dffr_apeg(ataf, jyro, d[0], apeg); // check edge
	assign #T_INV  aguz = !cpu_rd;
	assign #T_INV  byma = !ff24;
	assign #T_NOR  befu = !(aguz || byma);
	assign #T_INV  adak = !befu;
	assign #T_NAND bosu = !(ff24 && apu_wr);
	assign #T_INV  baxy = !bosu;
	assign #T_INV  bubu = !baxy;
	assign #T_INV  bowe = !bosu;
	assign #T_INV  ataf = !bowe;
	assign #T_TRI  atum = !adak ? bedu : 1'bz; /* takes !q output of dff */
	assign #T_TRI  bocy = !adak ? cozu : 1'bz; /* takes !q output of dff */
	assign #T_TRI  arux = !adak ? bumo : 1'bz; /* takes !q output of dff */
	assign #T_TRI  amad = !adak ? byre : 1'bz; /* takes !q output of dff */
	assign #T_TRI  axem = !adak ? apos : 1'bz; /* takes !q output of dff */
	assign #T_TRI  avud = !adak ? ager : 1'bz; /* takes !q output of dff */
	assign #T_TRI  awed = !adak ? byga : 1'bz; /* takes !q output of dff */
	assign #T_TRI  akod = !adak ? apeg : 1'bz; /* takes !q output of dff */
	assign ncpu_rd = aguz;
	assign d[7]    = atum;
	assign d[6]    = bocy;
	assign d[5]    = arux;
	assign d[4]    = amad;
	assign d[3]    = axem;
	assign d[2]    = avud;
	assign d[1]    = awed;
	assign d[0]    = akod;

	wire gepa, hefa, gumu, bupo, bono, byfa;
	wire bogu, bafo, atuf, anev, bepu, befo, bume, bofa;
	wire capu, caga, boca, buzu, cere, cada, cavu, cudu;
	dffr dffr_bogu(bono, jyro, d[1], bogu); // check edge
	dffr dffr_bafo(bono, jyro, d[2], bafo); // check edge
	dffr dffr_atuf(bono, jyro, d[3], atuf); // check edge
	dffr dffr_anev(bono, jyro, d[0], anev); // check edge
	dffr dffr_bepu(byfa, jyro, d[7], bepu); // check edge
	dffr dffr_befo(byfa, jyro, d[6], befo); // check edge
	dffr dffr_bume(byfa, jyro, d[4], bume); // check edge
	dffr dffr_bofa(byfa, jyro, d[5], bofa); // check edge
	assign #T_INV  gepa = !ff25;
	assign #T_NOR  hefa = !(ncpu_rd || gepa);
	assign #T_INV  gumu = !hefa;
	assign #T_NAND bupo = !(ff25 && apu_wr);
	assign #T_INV  bono = !bupo;
	assign #T_INV  byfa = !bupo;
	assign #T_TRI  capu = !gumu ? bogu : 1'bz; /* takes !q output of dff */
	assign #T_TRI  caga = !gumu ? bafo : 1'bz; /* takes !q output of dff */
	assign #T_TRI  boca = !gumu ? atuf : 1'bz; /* takes !q output of dff */
	assign #T_TRI  buzu = !gumu ? anev : 1'bz; /* takes !q output of dff */
	assign #T_TRI  cere = !gumu ? bepu : 1'bz; /* takes !q output of dff */
	assign #T_TRI  cada = !gumu ? befo : 1'bz; /* takes !q output of dff */
	assign #T_TRI  cavu = !gumu ? bume : 1'bz; /* takes !q output of dff */
	assign #T_TRI  cudu = !gumu ? bofa : 1'bz; /* takes !q output of dff */
	assign lmixer[1] = bogu;
	assign lmixer[2] = bafo;
	assign lmixer[3] = atuf;
	assign lmixer[0] = anev;
	assign rmixer[3] = bepu;
	assign rmixer[2] = befo;
	assign rmixer[0] = bume;
	assign rmixer[1] = bofa;
	assign d[1]      = capu;
	assign d[2]      = caga;
	assign d[3]      = boca;
	assign d[0]      = buzu;
	assign d[7]      = cere;
	assign d[6]      = cada;
	assign d[4]      = cavu;
	assign d[5]      = cudu;

	wire ceto, kazo, curu, dole, kamu, duru, fewa, coto, koge, efus, fate;
	assign #T_INV  ceto = !ncpu_rd;
	assign #T_INV  kazo = !ncpu_rd;
	assign #T_INV  curu = !ncpu_rd;
	assign #T_INV  gaxo = !ncpu_rd;
	assign #T_NAND dole = !(ff26 && ceto);
	assign #T_NAND kamu = !(ff26 && kazo);
	assign #T_NAND duru = !(ff26 && curu);
	assign #T_NAND fewa = !(ff26 && gaxo);
	assign #T_TRI  coto = !dole ? !nch1_active : 1'bz;
	assign #T_TRI  koge = !dole ? !nch4_active : 1'bz;
	assign #T_TRI  efus = !dole ? !nch2_active : 1'bz;
	assign #T_TRI  fate = !dole ? !nch3_active : 1'bz;
	assign d[0] = coto;
	assign d[3] = koge;
	assign d[1] = efus;
	assign d[2] = fate;

endmodule

module apu_decode(
		a,
		cpu_wr, cpu_rd,
		ff00wr, ff00rd, apu_wr, ff26, ff3x,
		ffxx, nffxx, anap, duce,
		nff1a_d7, nch1_amp_en, nch2_amp_en, nch4_amp_en, namp_en,
		ff10, ff11, ff12, ff13, ff14, ff16, ff17, ff18, ff19, ff1a,
		ff1b, ff1c, ff1d, ff1e, ff20, ff21, ff22, ff23, ff24, ff25
	);

	input wire [15:0] a;

	input wire cpu_wr, cpu_rd;

	output wire ff00wr, ff00rd, apu_wr, ff26, ff3x;
	input  wire ffxx, nffxx;
	output wire anap, duce;
	input  wire nff1a_d7, nch1_amp_en, nch2_amp_en, nch4_amp_en;
	output wire namp_en;

	output wire ff10, ff11, ff12, ff13, ff14, ff16, ff17, ff18, ff19, ff1a;
	output wire ff1b, ff1c, ff1d, ff1e, ff20, ff21, ff22, ff23, ff24, ff25;

	wire amus, byko, akug, atoz, acat;
	assign #T_NOR  amus = !(a[7] || a[4] || a[3] || a[2] || a[1] || a[0]);
	assign #T_AND  anap = amus && ffxx;
	assign #T_INV  byko = !a[5];
	assign #T_INV  akug = !a[6];
	assign #T_NAND atoz = !(byko && akug && cpu_wr && anap);
	assign #T_AND  acat = anap && cpu_rd && akug && byko;
	assign ff00wr = atoz;
	assign ff00rd = acat;

	wire boxy, awet, bezy, avun, asad, acom, baro, atup, ateg, buno, banu, cona, doxy, bafu, bogy, tace, nff1x;
	wire ff2x, nff2x;
	assign #T_INV  boxy = !a[5];
	assign #T_OR   awet = a[4] || boxy || a[6] || a[7];
	assign #T_OR   bezy = awet || nffxx;
	assign #T_INV  avun = !a[7];
	assign #T_INV  asad = !a[6];
	assign #T_NAND acom = !(avun && asad && a[5] && a[4]);
	assign #T_NOR  baro = !(acom || nffxx);
	assign #T_INV  atup = !a[4];
	assign #T_OR   ateg = atup || a[5] || a[6] || a[7];
	assign #T_NOR  buno = !(nffxx || ateg);
	assign #T_INV  banu = !buno;
	assign #T_INV  cona = !nff2x;
	assign #T_AND  doxy = cona && xxx6;
	assign #T_INV  bafu = !cpu_wr;
	assign #T_INV  bogy = !bafu;
	assign #T_AND  tace = nch1_amp_en && nch2_amp_en && nff1a_d7 && nch4_amp_en;
	assign nff2x   = bezy;
	assign ff3x    = baro;
	assign nff1x   = banu;
	assign ff2x    = cona;
	assign ff26    = doxy;
	assign apu_wr  = bogy;
	assign namp_en = tace;

	wire dyte, doso, afob, dupa, abub, deno, acol;
	wire dupo, datu, daza, dura, duvu, dofa, damy, dufe, duno, dewa, dejy, dona, dafy, emos;
	wire ekag, esot, egen, exat, emax, etuf, gany, dyva, cafy, covy, cora, dutu, ekez, edaf;
	wire cuge, caxe, covo, doza, danu, dara, feny, duja, dugo, emor, dusa, deco, gefo, xxx6;
	assign #T_INV  dyte = !a[0];
	assign #T_INV  doso = !dyte;
	assign #T_INV  afob = !a[1];
	assign #T_INV  dupa = !afob;
	assign #T_INV  abub = !a[2];
	assign #T_INV  deno = !abub;
	assign #T_INV  acol = !a[3];
	assign #T_INV  duce = !acol;
	assign #T_NAND dupo = !(acol && abub && afob && dyte);
	assign #T_NAND datu = !(dyte && afob && deno && acol);
	assign #T_NAND daza = !(acol && deno && dupa && dyte);
	assign #T_NAND dura = !(doso && afob && deno && acol);
	assign #T_NAND duvu = !(acol && deno && dupa && doso);
	assign #T_AND  dofa = acol && abub && dupa && dyte;
	assign #T_NAND damy = !(acol && abub && dupa && dyte);
	assign #T_NAND dufe = !(doso && dupa && abub && acol);
	assign #T_NAND duno = !(acol && abub && afob && doso);
	assign #T_NAND dewa = !(doso && afob && abub && acol);
	assign #T_NAND dejy = !(duce && abub && afob && doso);
	assign #T_NAND dona = !(dyte && afob && abub && acol);
	assign #T_NAND dafy = !(duce && abub && afob && dyte);
	assign #T_NAND emos = !(doso && afob && deno && duce);
	assign #T_AND  ekag = acol && deno && dupa && dyte;
	assign #T_NAND esot = !(acol && deno && afob && dyte);
	assign #T_NAND egen = !(dyte && dupa && deno && duce);
	assign #T_NAND exat = !(duce && abub && dupa && dyte);
	assign #T_NAND emax = !(doso && dupa && abub && duce);
	assign #T_NAND etuf = !(acol && abub && dupa && doso);
	assign #T_NAND gany = !(duce && deno && afob && dyte);
	assign #T_NOR  dyva = !(dupo || nff1x);
	assign #T_NOR  cafy = !(datu || nff2x);
	assign #T_NOR  covy = !(daza || nff1x);
	assign #T_NOR  cora = !(dura || nff2x);
	assign #T_NOR  dutu = !(duvu || nff1x);
	assign #T_AND  ekez = dofa && ff2x;
	assign #T_NOR  edaf = !(damy || nff1x);
	assign #T_NOR  cuge = !(dufe || nff2x);
	assign #T_NOR  caxe = !(duno || nff1x);
	assign #T_NOR  covo = !(dewa || nff2x);
	assign #T_NOR  doza = !(dejy || nff1x);
	assign #T_NOR  danu = !(dona || nff2x);
	assign #T_NOR  dara = !(dafy || nff1x);
	assign #T_NOR  feny = !(emos || nff1x);
	assign #T_NOR  duja = !(esot || nff1x);
	assign #T_NOR  dugo = !(egen || nff1x);
	assign #T_NOR  emor = !(exat || nff1x);
	assign #T_NOR  dusa = !(emax || nff1x);
	assign #T_NOR  deco = !(etuf || nff1x);
	assign #T_NOR  gefo = !(gany || nff1x);
	assign xxx6 = ekag;
	assign ff10 = dyva;
	assign ff24 = cafy;
	assign ff16 = covy;
	assign ff25 = cora;
	assign ff17 = dutu;
	assign ff22 = ekez;
	assign ff12 = edaf;
	assign ff23 = cuge;
	assign ff11 = caxe;
	assign ff21 = covo;
	assign ff19 = doza;
	assign ff20 = danu;
	assign ff18 = dara;
	assign ff1d = feny;
	assign ff14 = duja;
	assign ff1e = dugo;
	assign ff1a = emor;
	assign ff1b = dusa;
	assign ff13 = deco;
	assign ff1c = gefo;

endmodule

module vram_ifc(
		a, ma, ma_out,
		md, md_in, md_out, md_a,
		d, d_in, d_a,
		oam_a_d, oam_b_d,
		moe_in, mwr_in, mcs_in, moe_a, moe_d, mwr_a, mwr_d, mcs_a, mcs_d, md_b,
		nt1_t2, dma_run, mopa_phi, nfexxffxx, nreset6, cpu_rd_sync, vram_to_oam, dma_addr_ext, ff40_d4,
		roru, lula, bedo, saro, tacu, tuvo, acyl, xyso, texo, abuz, afas, texy, myma, lena, xymu, leko,
		xuha, vyno, vujo, vymu, neta, pore, potu, npyju, npowy, npoju, npulo, npoxa, npyzo, npozo, nrawu,
		cota, wuko
	);

	input wire [15:0] a;

	inout  wire [12:0] ma;
	output wire [12:0] ma_out;

	inout  wire [7:0] d;
	input  wire [7:0] d_in;
	output wire [7:0] d_a;

	inout  wire [7:0] md;
	input  wire [7:0] md_in;
	output wire [7:0] md_out, md_a;

	output wire [7:0] oam_a_d, oam_b_d;

	input  wire moe_in, mwr_in, mcs_in;
	output wire moe_a, moe_d, mwr_a, mwr_d, mcs_a, mcs_d, md_b;

	input wire nt1_t2, dma_run, mopa_phi, nfexxffxx, nreset6, cpu_rd_sync, vram_to_oam, dma_addr_ext, ff40_d4;

	input  wire roru, lula, bedo, saro, tacu, tuvo, acyl, xyso, texo, abuz, afas, texy, myma, lena, xymu, leko;
	input  wire xuha, vyno, vujo, vymu, neta, pore, potu, npyju, npowy, npoju, npulo, npoxa, npyzo, npozo, nrawu;
	output wire cota, wuko;

	wire reho, pony, ruma, pedu, ruky, nuva, vode, tago, vova, tujy, mume, luby, mewy;
	wire lefa, mysa, lalo, mepa, loly, mavu, luvo, myre, laca, masa, lozu, myfu, lexe;
	assign #T_INV  reho = !ma[12];
	assign #T_INV  ruma = !ma[11];
	assign #T_INV  ruky = !ma[10];
	assign #T_INV  vode = !ma[9];
	assign #T_INV  vova = !ma[8];
	assign #T_INV  mume = !ma[7];
	assign #T_INV  mewy = !ma[6];
	assign #T_INV  mysa = !ma[5];
	assign #T_INV  mepa = !ma[4];
	assign #T_INV  mavu = !ma[3];
	assign #T_INV  myre = !ma[2];
	assign #T_INV  masa = !ma[1];
	assign #T_INV  myfu = !ma[0];
	assign #T_INV  pony = !reho;
	assign #T_INV  pedu = !ruma;
	assign #T_INV  nuva = !ruky;
	assign #T_INV  tago = !vode;
	assign #T_INV  tujy = !vova;
	assign #T_INV  luby = !mume;
	assign #T_INV  lefa = !mewy;
	assign #T_INV  lalo = !mysa;
	assign #T_INV  loly = !mepa;
	assign #T_INV  luvo = !mavu;
	assign #T_INV  laca = !myre;
	assign #T_INV  lozu = !masa;
	assign #T_INV  lexe = !myfu;
	assign ma_out[12] = pony;
	assign ma_out[11] = pedu;
	assign ma_out[10] = nuva;
	assign ma_out[9]  = tago;
	assign ma_out[8]  = tujy;
	assign ma_out[7]  = luby;
	assign ma_out[6]  = lefa;
	assign ma_out[5]  = lalo;
	assign ma_out[4]  = loly;
	assign ma_out[3]  = luvo;
	assign ma_out[2]  = laca;
	assign ma_out[1]  = lozu;
	assign ma_out[0]  = lexe;

	wire ryvo, rera, raby, rory, ruja, ravu, rafy, ruxa;
	assign #T_NAND ryvo = !(d[5] && lula);
	assign #T_NAND rera = !(d[3] && lula);
	assign #T_NAND raby = !(d[2] && lula);
	assign #T_NAND rory = !(d[4] && lula);
	assign #T_NAND ruja = !(d[1] && lula);
	assign #T_NAND ravu = !(d[7] && lula);
	assign #T_NAND rafy = !(d[6] && lula);
	assign #T_NAND ruxa = !(d[0] && lula);
	assign d_a[5] = ryvo;
	assign d_a[3] = rera;
	assign d_a[2] = raby;
	assign d_a[4] = rory;
	assign d_a[1] = ruja;
	assign d_a[7] = ravu;
	assign d_a[6] = rafy;
	assign d_a[0] = ruxa;

	wire cufe, vape, aver, xujy, bycu;
	assign #T_NAO  cufe = !((saro && dma_run) || mopa_phi);
	assign #T_AND  vape = tacu && tuvo;
	assign #T_AND  aver = acyl && xyso;
	assign #T_INV  xujy = !vape;
	assign #T_NOR  bycu = !(cufe || xujy || aver);
	assign #T_INV  cota = !bycu;

	wire syro, tefa, sose, tuca, tuja, tegu, tavy, sycy, soto, tuto, sudo, tefy, sale, tyjy, tole;
	dffr dffr_soto(sycy, nreset6, !soto, soto); // check edge
	assign #T_INV  syro = !nfexxffxx;
	assign #T_NOR  tefa = !(syro || texo);
	assign #T_AND  sose = a[15] && tefa;
	assign #T_AND  tuca = sose && abuz;
	assign #T_AND  tuja = sose && cpu_rd_sync;
	assign #T_NAND tegu = !(sose && afas);
	assign #T_INV  tavy = !moe_in;
	assign #T_INV  sycy = !nt1_t2;
	assign #T_AND  tuto = nt1_t2 && !soto;
	assign #T_INV  sudo = !mwr_in;
	assign #T_INV  tefy = !mcs_in;
	assign #T_MUX  sale = tuto ? tavy : tegu;
	assign #T_MUX  tyjy = tuto ? sudo : tuja;
	assign #T_MUX  tole = tuto ? tefy : tuca;

	wire soho, rawa, raco, rylu, racu, apam, ruvy, sohy, sutu, sere, sazo, ropy, ryje, revo, rela, rocy;
	wire rena, rahu, rofa, rute, sema, sofy, taxy, sewo, tode, saha, refo, ragu, sysy, sety, soky;
	assign #T_AND  soho = tacu && texy;
	assign #T_INV  rawa = !soho;
	assign #T_NAND rylu = !(sale && ropy);
	assign #T_INV  apam = !vram_to_oam;
	assign #T_AND  racu = rylu && rawa && myma && apam;
	assign #T_INV  raco = !tuto;
	assign #T_INV  ruvy = !sale;
	assign #T_NOR  sutu = !(lena || vram_to_oam || texy || sere);
	assign #T_NAND sohy = !(tyjy && sere);
	assign #T_INV  ropy = !xymu;
	assign #T_AND  sere = tole && ropy;
	assign #T_AND  sazo = ruvy && sere;
	assign #T_INV  ryje = !sazo;
	assign #T_INV  revo = !ryje;
	assign #T_OR   rela = revo || sazo;
	assign #T_INV  rena = !rela;
	assign #T_INV  rofa = !rena;
	assign #T_AND  rocy = sazo && revo;
	assign #T_INV  rahu = !rocy;
	assign #T_OR   rute = tuto || raco;
	assign #T_AND  sema = racu && raco;
	assign #T_OR   sofy = tuto || sohy;
	assign #T_AND  taxy = sohy && raco;
	assign #T_OR   sewo = tuto || sutu;
	assign #T_AND  tode = sutu && raco;
	assign #T_INV  saha = !rute;
	assign #T_INV  refo = !sema;
	assign #T_INV  ragu = !sofy;
	assign #T_INV  sysy = !taxy;
	assign #T_INV  sety = !sewo;
	assign #T_INV  soky = !tode;
	assign moe_d = saha;
	assign moe_a = refo;
	assign mwr_d = ragu;
	assign mwr_a = sysy;
	assign mcs_d = sety;
	assign mcs_a = soky;
	assign md_b = rofa;

	wire raku, roce, remo, ropu, reta, rydo, rody, reba;
	assign #T_TRI  raku = rena ? !md_in[7] : 1'bz;
	assign #T_TRI  roce = rena ? !md_in[4] : 1'bz;
	assign #T_TRI  remo = rena ? !md_in[3] : 1'bz;
	assign #T_TRI  ropu = rena ? !md_in[5] : 1'bz;
	assign #T_TRI  reta = rena ? !md_in[6] : 1'bz;
	assign #T_TRI  rydo = rena ? !md_in[2] : 1'bz;
	assign #T_TRI  rody = rena ? !md_in[0] : 1'bz;
	assign #T_TRI  reba = rena ? !md_in[1] : 1'bz;
	assign md[7] = raku;
	assign md[4] = roce;
	assign md[3] = remo;
	assign md[5] = ropu;
	assign md[6] = reta;
	assign md[2] = rydo;
	assign md[0] = rody;
	assign md[1] = reba;

	wire runy, tuso, sole, tahy, tesu, taxo, tovu, tazu, tewa, sosa, sedu;
	assign         runy = 1'b1;
	assign #T_NOR  tuso = !(nt1_t2 || bedo);
	assign #T_INV  sole = !tuso;
	assign #T_TRI  tahy = !runy ? !sole : 1'bz; // check enable input polarity
	assign #T_TRI  tesu = !runy ? !sole : 1'bz; // check enable input polarity
	assign #T_TRI  taxo = !runy ? !sole : 1'bz; // check enable input polarity
	assign #T_TRI  tovu = !runy ? !sole : 1'bz; // check enable input polarity
	assign #T_TRI  tazu = !runy ? !sole : 1'bz; // check enable input polarity
	assign #T_TRI  tewa = !runy ? !sole : 1'bz; // check enable input polarity
	assign #T_TRI  sosa = !runy ? !sole : 1'bz; // check enable input polarity
	assign #T_TRI  sedu = !runy ? !sole : 1'bz; // check enable input polarity
	assign d[4] = tahy;
	assign d[5] = tesu;
	assign d[3] = taxo;
	assign d[0] = tovu;
	assign d[6] = tazu;
	assign d[7] = tewa;
	assign d[1] = sosa;
	assign d[2] = sedu;

	wire xane, xedu, xeca, xybo, rysu, ruse, rumo, xyne, xoba, xody, ryna, rese, xaky, xopo, xuxu;
	assign #T_NOR  xane = !(vram_to_oam || xymu);
	assign #T_INV  xedu = !xane;
	assign #T_TRI  xeca = !xedu ? !a[4]  : 1'bz;
	assign #T_TRI  xybo = !xedu ? !a[7]  : 1'bz;
	assign #T_TRI  rysu = !xedu ? !a[8]  : 1'bz;
	assign #T_TRI  ruse = !xedu ? !a[10] : 1'bz;
	assign #T_TRI  rumo = !xedu ? !a[12] : 1'bz;
	assign #T_TRI  xyne = !xedu ? !a[2]  : 1'bz;
	assign #T_TRI  xoba = !xedu ? !a[5]  : 1'bz;
	assign #T_TRI  xody = !xedu ? !a[3]  : 1'bz;
	assign #T_TRI  ryna = !xedu ? !a[11] : 1'bz;
	assign #T_TRI  rese = !xedu ? !a[9]  : 1'bz;
	assign #T_TRI  xaky = !xedu ? !a[0]  : 1'bz;
	assign #T_TRI  xopo = !xedu ? !a[6]  : 1'bz;
	assign #T_TRI  xuxu = !xedu ? !a[1]  : 1'bz;
	assign ma[4]  = xeca;
	assign ma[7]  = xybo;
	assign ma[8]  = rysu;
	assign ma[10] = ruse;
	assign ma[12] = rumo;
	assign ma[2]  = xyne;
	assign ma[5]  = xoba;
	assign ma[3]  = xody;
	assign ma[11] = ryna;
	assign ma[9]  = rese;
	assign ma[0]  = xaky;
	assign ma[6]  = xopo;
	assign ma[1]  = xuxu;

	wire lyra, ryba, ruzy, rome, tehe, soca, ratu, tovo, saza;
	wire ropa, sywa, sugu, tute, temy, sajo, tuty, tawo;
	assign #T_NAND lyra = !(nt1_t2 && roru);
	assign #T_INV  ryba = !d_in[7];
	assign #T_INV  ruzy = !d_in[1];
	assign #T_INV  rome = !d_in[2];
	assign #T_INV  tehe = !d_in[4];
	assign #T_INV  soca = !d_in[6];
	assign #T_INV  ratu = !d_in[5];
	assign #T_INV  tovo = !d_in[0];
	assign #T_INV  saza = !d_in[3];
	assign #T_TRI  ropa = !lyra ? !ryba : 1'bz; // check enable input polarity
	assign #T_TRI  sywa = !lyra ? !ruzy : 1'bz; // check enable input polarity
	assign #T_TRI  sugu = !lyra ? !rome : 1'bz; // check enable input polarity
	assign #T_TRI  tute = !lyra ? !tehe : 1'bz; // check enable input polarity
	assign #T_TRI  temy = !lyra ? !soca : 1'bz; // check enable input polarity
	assign #T_TRI  sajo = !lyra ? !ratu : 1'bz; // check enable input polarity
	assign #T_TRI  tuty = !lyra ? !tovo : 1'bz; // check enable input polarity
	assign #T_TRI  tawo = !lyra ? !saza : 1'bz; // check enable input polarity
	assign d[7] = ropa;
	assign d[1] = sywa;
	assign d[2] = sugu;
	assign d[4] = tute;
	assign d[6] = temy;
	assign d[5] = sajo;
	assign d[0] = tuty;
	assign d[3] = tawo;

	wire rove, sefa, suna, sumo, suke, samo, sogo, sazu, sefu, rege, rada, ryro, ryze, reku, ryky, revu, razo;
	assign #T_INV  rove = !rahu;
	assign #T_AND  sefa = md[0] && rove;
	assign #T_AND  suna = md[3] && rove;
	assign #T_AND  sumo = md[4] && rove;
	assign #T_AND  suke = md[7] && rove;
	assign #T_AND  samo = md[6] && rove;
	assign #T_AND  sogo = md[1] && rove;
	assign #T_AND  sazu = md[5] && rove;
	assign #T_AND  sefu = md[2] && rove;
	assign #T_INV  rege = !sefa;
	assign #T_INV  rada = !suna;
	assign #T_INV  ryro = !sumo;
	assign #T_INV  ryze = !suke;
	assign #T_INV  reku = !samo;
	assign #T_INV  ryky = !sogo;
	assign #T_INV  revu = !sazu;
	assign #T_INV  razo = !sefu;
	assign md_a[0] = rege;
	assign md_a[3] = rada;
	assign md_a[4] = ryro;
	assign md_a[7] = ryze;
	assign md_a[6] = reku;
	assign md_a[1] = ryky;
	assign md_a[5] = revu;
	assign md_a[2] = razo;

	wire cede, syzo, tune, sera, sysa, tube, sugy, ralo, tenu;
	wire bape, bypy, bomo, bubo, basa, betu, buma, baxu, basy, byny, bupy, buhu, wasa, wejo, cako, cyme;
	assign #T_INV  cede = !dma_addr_ext;
	assign #T_INV  syzo = !d_in[7];
	assign #T_INV  tune = !d_in[1];
	assign #T_INV  sera = !d_in[2];
	assign #T_INV  sysa = !d_in[4];
	assign #T_INV  tube = !d_in[6];
	assign #T_INV  sugy = !d_in[5];
	assign #T_INV  ralo = !d_in[0];
	assign #T_INV  tenu = !d_in[3];
	assign #T_TRI  bape = !cede ? !syzo : 1'bz;
	assign #T_TRI  bypy = !cede ? !syzo : 1'bz;
	assign #T_TRI  bomo = !cede ? !tune : 1'bz;
	assign #T_TRI  bubo = !cede ? !tune : 1'bz;
	assign #T_TRI  basa = !cede ? !sera : 1'bz;
	assign #T_TRI  betu = !cede ? !sera : 1'bz;
	assign #T_TRI  buma = !cede ? !sysa : 1'bz;
	assign #T_TRI  baxu = !cede ? !sysa : 1'bz;
	assign #T_TRI  basy = !cede ? !tube : 1'bz;
	assign #T_TRI  byny = !cede ? !tube : 1'bz;
	assign #T_TRI  bupy = !cede ? !sugy : 1'bz;
	assign #T_TRI  buhu = !cede ? !sugy : 1'bz;
	assign #T_TRI  wasa = !cede ? !ralo : 1'bz;
	assign #T_TRI  wejo = !cede ? !ralo : 1'bz;
	assign #T_TRI  cako = !cede ? !tenu : 1'bz;
	assign #T_TRI  cyme = !cede ? !tenu : 1'bz;
	assign oam_b_d[7] = bape;
	assign oam_a_d[7] = bypy;
	assign oam_b_d[1] = bomo;
	assign oam_a_d[1] = bubo;
	assign oam_a_d[2] = basa;
	assign oam_b_d[2] = betu;
	assign oam_b_d[4] = buma;
	assign oam_a_d[4] = baxu;
	assign oam_b_d[6] = basy;
	assign oam_a_d[6] = byny;
	assign oam_a_d[5] = bupy;
	assign oam_b_d[5] = buhu;
	assign oam_a_d[0] = wasa;
	assign oam_b_d[0] = wejo;
	assign oam_b_d[3] = cako;
	assign oam_a_d[3] = cyme;

	wire tyvy, seby, roro, rery, rona, runa, runo, same, sana, rabo, rexu, ruga, rybu, rota, raju, toku, tyja, rupy;
	assign #T_NAND tyvy = !(sere && leko);
	assign #T_INV  seby = !tyvy;
	assign #T_INV  roro = !md[5];
	assign #T_INV  rery = !md[0];
	assign #T_INV  rona = !md[2];
	assign #T_INV  runa = !md[1];
	assign #T_INV  runo = !md[3];
	assign #T_INV  same = !md[7];
	assign #T_INV  sana = !md[4];
	assign #T_INV  rabo = !md[6];
	assign #T_TRI  rexu = seby ? !roro : 1'bz;
	assign #T_TRI  ruga = seby ? !rery : 1'bz;
	assign #T_TRI  rybu = seby ? !rona : 1'bz;
	assign #T_TRI  rota = seby ? !runa : 1'bz;
	assign #T_TRI  raju = seby ? !runo : 1'bz;
	assign #T_TRI  toku = seby ? !same : 1'bz;
	assign #T_TRI  tyja = seby ? !sana : 1'bz;
	assign #T_TRI  rupy = seby ? !rabo : 1'bz;
	assign d[5] = rexu;
	assign d[0] = ruga;
	assign d[2] = rybu;
	assign d[1] = rota;
	assign d[3] = raju;
	assign d[7] = toku;
	assign d[4] = tyja;
	assign d[6] = rupy;

	wire xonu, wudo, wawe, wolu, xucy, xeze;
	assign #T_TRI  xonu = !xucy ? !xuha : 1'bz;
	assign #T_TRI  wudo = !xucy ? !vyno : 1'bz;
	assign #T_TRI  wawe = !xucy ? !vujo : 1'bz;
	assign #T_TRI  wolu = !xucy ? !vymu : 1'bz;
	assign #T_NAND xucy = !(neta && pore);
	assign #T_AND  xeze = potu && pore;
	assign #T_INV  wuko = !xeze;

	wire teme, tewu, tygo, sote, seke, rujo, tofa, suza;
	wire synu, syma, roko, sybu, sako, sejy, sedo, sawu;
	wire rura, ruly, rare, rodu, rube, rumu, ryty, rady;
	assign #T_TRI  teme = !rahu ? !d[0] : 1'bz; // check enable input polarity
	assign #T_TRI  tewu = !rahu ? !d[1] : 1'bz; // check enable input polarity
	assign #T_TRI  tygo = !rahu ? !d[2] : 1'bz; // check enable input polarity
	assign #T_TRI  sote = !rahu ? !d[3] : 1'bz; // check enable input polarity
	assign #T_TRI  seke = !rahu ? !d[4] : 1'bz; // check enable input polarity
	assign #T_TRI  rujo = !rahu ? !d[5] : 1'bz; // check enable input polarity
	assign #T_TRI  tofa = !rahu ? !d[6] : 1'bz; // check enable input polarity
	assign #T_TRI  suza = !rahu ? !d[7] : 1'bz; // check enable input polarity
	assign #T_OR   synu = rahu || md[0];
	assign #T_OR   syma = rahu || md[1];
	assign #T_OR   roko = rahu || md[2];
	assign #T_OR   sybu = rahu || md[3];
	assign #T_OR   sako = rahu || md[4];
	assign #T_OR   sejy = rahu || md[5];
	assign #T_OR   sedo = rahu || md[6];
	assign #T_OR   sawu = rahu || md[7];
	assign #T_INV  rura = !synu;
	assign #T_INV  ruly = !syma;
	assign #T_INV  rare = !roko;
	assign #T_INV  rodu = !sybu;
	assign #T_INV  rube = !sako;
	assign #T_INV  rumu = !sejy;
	assign #T_INV  ryty = !sedo;
	assign #T_INV  rady = !sawu;
	assign md[0] = teme;
	assign md[1] = tewu;
	assign md[2] = tygo;
	assign md[3] = sote;
	assign md[4] = seke;
	assign md[5] = rujo;
	assign md[6] = tofa;
	assign md[7] = suza;
	assign md_out[0] = rura;
	assign md_out[1] = ruly;
	assign md_out[2] = rare;
	assign md_out[3] = rodu;
	assign md_out[4] = rube;
	assign md_out[5] = rumu;
	assign md_out[6] = ryty;
	assign md_out[7] = rady;

	wire vuza, vury, tobo, suvo, reso, roha, rusa, vejy, sezu, vapy;
	assign #T_NOR  vuza = !(ff40_d4 || npyju);
	assign #T_TRI  vury = neta ? !vuza  : 1'bz;
	assign #T_TRI  tobo = neta ? !npyju : 1'bz;
	assign #T_TRI  suvo = neta ? !npowy : 1'bz;
	assign #T_TRI  reso = neta ? !npoju : 1'bz;
	assign #T_TRI  roha = neta ? !npulo : 1'bz;
	assign #T_TRI  rusa = neta ? !npoxa : 1'bz;
	assign #T_TRI  vejy = neta ? !npyzo : 1'bz;
	assign #T_TRI  sezu = neta ? !npozo : 1'bz;
	assign #T_TRI  vapy = neta ? !nrawu : 1'bz;
	assign ma[12] = vury;
	assign ma[11] = tobo;
	assign ma[10] = suvo;
	assign ma[9]  = reso;
	assign ma[8]  = roha;
	assign ma[7]  = rusa;
	assign ma[6]  = vejy;
	assign ma[5]  = sezu;
	assign ma[4]  = vapy;

endmodule

module dffr(clk, nreset, d, q);

	parameter INITIAL_Q = 2;

	input  wire clk, nreset, d;
	output wire q;

	reg ff;

	initial if (INITIAL_Q != 0 && INITIAL_Q != 1) ff = $random; else ff = INITIAL_Q;

	always @(posedge clk or negedge nreset) begin
		if (nreset)
			ff <= (d === 1'bx) ? $random : d;
		else
			ff <= 0;
	end

	assign #T_DFFR q = ff;

endmodule

module dff(clk, d, q);

	parameter INITIAL_Q = 2;

	input  wire clk, d;
	output wire q;

	reg ff;

	initial if (INITIAL_Q != 0 && INITIAL_Q != 1) ff = $random; else ff = INITIAL_Q;

	always @(posedge clk) begin
		ff <= (d === 1'bx) ? $random : d;
	end

	assign #T_DFF q = ff;

endmodule

module latch(c, d, q);

	input  wire c, d;
	output wire q;

	assign #T_LATCH q = c ? d : q;

endmodule
