`default_nettype none

module sm83_nor2_pch_in1_dec3 #(
		parameter real L_in1 = 27,
		parameter real L_y   = 45
	) (
		input     logic pch_n, in2,
		inout tri logic in1,
		output    logic y
	);

	import sm83_timing::*;

	assign y = !(in1 | in2);

	localparam realtime T_rise_buf = tpd_elmore(L_in1, R_pmos_ohm(8*L_unit));
	localparam realtime T_Z_buf    = tpd_z(T_rise_buf);
	bufif0 (strong1, highz0) #(T_rise_buf, 0, T_Z_buf) (in1, '1, pch_n);

	specify
		specparam T_rise_y = tpd_elmore(L_y, R_pmos_ohm(17*L_unit) * 2);
		specparam T_fall_y = tpd_elmore(L_y, R_nmos_ohm( 8*L_unit));

		(in1, in2 *> y) = (T_rise_y, T_fall_y);
	endspecify

endmodule

`default_nettype wire
