`default_nettype none

module sprite_control(
		inout tri logic [7:0]  d,
		input logic     [7:0]  oam_b_nd, v,
		inout tri logic [12:0] nma,

		input logic clk1, clk2, clk3, clk4, clk5, reset_video, nreset_video, oam_b_cpu_nrd,

		input logic ff40_d1, ff40_d2,

		input  logic nxymu, ynaz, ykok, zure, ywos, ekes, cehu, ewam, cyvy, zako, xeba,
		input  logic ylev, ytub, feha, dama, cyco, daje, ydot, ywap, fyma, cogy, byva,
		input  logic cota, nyzos, sela, xyvo, anom, feto, seca, nbaxo, azyb,
		input  logic wenu, cucu, cuca, cega, besu,
		output logic fepo, fado, deny, gugy, xyme, gygy, gowo, gyma, fame, dydo, furo,
		output logic wuty, dosy, wuzo, gafy, xaho, ejad, wunu, wupa, gamy, doku, dyna,
		output logic texy, dege, daby, dabu, gysa, wuvu_nq, xupy, abez, xoce, catu, xyso,
		output logic buza, avap, tyfo_nq, tuvo, tacu, xefy, xono, xado, puco,
		output logic cacu, buzy, fuke, zape, wuse, zuru, fefo, gecy, wabe,
		output logic feka, xyha, yfag, cexu, akol, bymy, fuxu, enob, geny,
		output logic weme, wufa, faka, cyla, dymo, bucy, wofo, wylu, ewot,
		output logic asys, ahof, byvy
	);

	logic byjo, azem, aror, xage, yloz, dego, dydu, ydug, ygem, efyl, dyka, ybez, egom;
	logic fefy, fove, wefu, geze, guva, gaja, fuma, enut, gupo, gede, emol, webo, wuto;
	logic gyfy, wuna, xyla, gono, gaba, weja, gega, wase, wyla, xoja, gyte, favo, gutu;
	logic geke, gyga, foxa, guze;
	logic dyba, fono, exuq, wapo, womy, wafy, xudy, gota, egav, cedy, eboj;
	logic dubu, goro, guky, wacy, feve, wohu, gake, foko, efev, dywe;
	dffr_bp dffr_fono(wuty, byva, guze, fono);
	dffr_bp dffr_exuq(wuty, byva, foxa, exuq);
	dffr_bp dffr_wapo(wuty, byva, gutu, wapo);
	dffr_bp dffr_womy(wuty, byva, xoja, womy);
	dffr_bp dffr_wafy(wuty, byva, gega, wafy);
	dffr_bp dffr_xudy(wuty, byva, gono, xudy);
	dffr_bp dffr_gota(wuty, byva, gyfy, gota);
	dffr_bp dffr_egav(wuty, byva, emol, egav);
	dffr_bp dffr_cedy(wuty, byva, enut, cedy);
	dffr_bp dffr_eboj(wuty, byva, guva, eboj);
	assign  byjo = !ceha;
	assign  azem = byjo && nxymu;
	assign  aror = azem && ff40_d1;
	assign xage = !(aror && ynaz && ykok);
	assign yloz = !(aror && zure && ywos);
	assign dego = !(aror && ekes && cehu);
	assign dydu = !(aror && ewam && cyvy);
	assign ydug = !(aror && zako && xeba);
	assign ygem = !(aror && ylev && ytub);
	assign efyl = !(aror && feha && dama);
	assign dyka = !(aror && cyco && daje);
	assign ybez = !(aror && ydot && ywap);
	assign egom = !(aror && fyma && cogy);
	assign fefy = !(xage && yloz && dego && dydu && ydug);
	assign fove = !(ygem && efyl && dyka && ybez && egom);
	assign   fepo = fefy || fove;
	assign  wefu = !ydug;
	assign   geze = wefu || '0;
	assign  guva = !(ydug || '0);
	assign  gaja = !dydu;
	assign   fuma = gaja || geze;
	assign  enut = !(dydu || geze);
	assign  gupo = !dego;
	assign   gede = gupo || fuma;
	assign  emol = !(dego || fuma);
	assign  webo = !yloz;
	assign   wuto = webo || gede;
	assign  gyfy = !(yloz || gede);
	assign  wuna = !xage;
	assign   xyla = wuna || wuto;
	assign  gono = !(xage || wuto);
	assign  gaba = !egom;
	assign   weja = gaba || xyla;
	assign  gega = !(egom || xyla);
	assign  wase = !ybez;
	assign   wyla = wase || weja;
	assign  xoja = !(ybez || weja);
	assign  gyte = !dyka;
	assign   favo = gyte || wyla;
	assign  gutu = !(dyka || wyla);
	assign  geke = !efyl;
	assign   gyga = geke || favo;
	assign  foxa = !(efyl || favo);
	assign  guze = !(ygem || gyga);
	assign  fado = !guze;
	assign  deny = !foxa;
	assign  gugy = !gutu;
	assign  xyme = !xoja;
	assign  gygy = !gega;
	assign  gowo = !gono;
	assign  gyma = !gyfy;
	assign  fame = !emol;
	assign  dydo = !enut;
	assign  furo = !guva;
	assign  dyba = !byva;
	assign   dubu = dyba || fono;
	assign   goro = dyba || exuq;
	assign   guky = dyba || wapo;
	assign   wacy = dyba || womy;
	assign   feve = dyba || wafy;
	assign   wohu = dyba || xudy;
	assign   gake = dyba || gota;
	assign   foko = dyba || egav;
	assign   efev = dyba || cedy;
	assign   dywe = dyba || eboj;
	assign  dosy = !dubu;
	assign  wuzo = !goro;
	assign  gafy = !guky;
	assign  xaho = !wacy;
	assign  ejad = !feve;
	assign  wunu = !wohu;
	assign  wupa = !gake;
	assign  gamy = !foko;
	assign  doku = !efev;
	assign  dyna = !dywe;

	logic yceb, zuca, WONE, zaxe, xafu, yses, zeca, ydyv;
	logic xele, ypon, xuvo, zysa, yweg, xabu, ytux, yfap;
	logic ywok, xegu, yjex, xyju, ybog, wyso, xote, yzab, xuso;
	logic abon, fugy, gavo, wyga, wune, gotu, gegu, xehe;
	logic ebos, dasa, fuky, fuve, fepu, fofa, femo, gusu;
	logic eruc, enef, feco, gyky, gopu, fuwa, goju, wuhu;
	logic eruc_c, enef_c, feco_c, gyky_c, gopu_c, fuwa_c, goju_c, wuhu_c;
	logic gace, guvu, gyda, gewy, govu, wota, gese, spr_match;
	logic tobu, vonu, wuky, wago, cyvu, bore, buvy, xuqu;
	logic baxe, aras, agag, abem, dyso, fufo, gejy, famu;
	dffr_bp dffr_tobu(clk5, nxymu, tuly, tobu);
	dffr_bp dffr_vonu(clk5, nxymu, tobu, vonu);
	dlatch_a latch_xegu(!ywok, yceb, xegu);
	dlatch_a latch_yjex(!ywok, zuca, yjex);
	dlatch_a latch_xyju(!ywok, WONE, xyju);
	dlatch_a latch_ybog(!ywok, zaxe, ybog);
	dlatch_a latch_wyso(!ywok, xafu, wyso);
	dlatch_a latch_xote(!ywok, yses, xote);
	dlatch_a latch_yzab(!ywok, zeca, yzab);
	dlatch_a latch_xuso(!ywok, ydyv, xuso);
	dlatch_b latch_yceb(clk3, oam_b_nd[1], yceb);
	dlatch_b latch_zuca(clk3, oam_b_nd[2], zuca);
	dlatch_b latch_wone(clk3, oam_b_nd[3], WONE);
	dlatch_b latch_zaxe(clk3, oam_b_nd[4], zaxe);
	dlatch_b latch_xafu(clk3, oam_b_nd[5], xafu);
	dlatch_b latch_yses(clk3, oam_b_nd[6], yses);
	dlatch_b latch_zeca(clk3, oam_b_nd[7], zeca);
	dlatch_b latch_ydyv(clk3, oam_b_nd[0], ydyv);
	assign xele = !oam_b_cpu_nrd ? !yceb : 'z;
	assign ypon = !oam_b_cpu_nrd ? !zuca : 'z;
	assign xuvo = !oam_b_cpu_nrd ? !WONE : 'z;
	assign zysa = !oam_b_cpu_nrd ? !zaxe : 'z;
	assign yweg = !oam_b_cpu_nrd ? !xafu : 'z;
	assign xabu = !oam_b_cpu_nrd ? !yses : 'z;
	assign ytux = !oam_b_cpu_nrd ? !zeca : 'z;
	assign yfap = !oam_b_cpu_nrd ? !ydyv : 'z;
	assign  ywok = !cota;
	assign  abon = !texy;
	assign  fugy = !abon ? !(!xegu) : 'z;
	assign  gavo = !abon ? !(!yjex) : 'z;
	assign  wyga = !abon ? !(!xyju) : 'z;
	assign  wune = !abon ? !(!ybog) : 'z;
	assign  gotu = !abon ? !(!wyso) : 'z;
	assign  gegu = !abon ? !(!xote) : 'z;
	assign  xehe = !abon ? !(!yzab) : 'z;
	assign  ebos = !v[0];
	assign  dasa = !v[1];
	assign  fuky = !v[2];
	assign  fuve = !v[3];
	assign  fepu = !v[4];
	assign  fofa = !v[5];
	assign  femo = !v[6];
	assign  gusu = !v[7];
	assign  { eruc_c, eruc } = ebos + !xuso + '0;
	assign  { enef_c, enef } = dasa + !xegu + eruc_c;
	assign  { feco_c, feco } = fuky + !yjex + enef_c;
	assign  { gyky_c, gyky } = fuve + !xyju + feco_c;
	assign  { gopu_c, gopu } = fepu + !ybog + gyky_c;
	assign  { fuwa_c, fuwa } = fofa + !wyso + gopu_c;
	assign  { goju_c, goju } = femo + !xote + fuwa_c;
	assign  { wuhu_c, wuhu } = gusu + !yzab + goju_c;
	assign  dege = !eruc;
	assign  daby = !enef;
	assign  dabu = !feco;
	assign  gysa = !gyky;
	assign  gace = !gopu;
	assign  guvu = !fuwa;
	assign  gyda = !goju;
	assign  gewy = !wuhu;
	assign   govu = ff40_d2 || gyky;
	assign wota = !(gace && guvu && gyda && gewy && wuhu_c && govu);
	assign  gese = !wota;
	assign  wuky = !nyzos;
	assign  wago = wuky != wenu;
	assign  cyvu = wuky != cucu;
	assign  bore = wuky != cuca;
	assign  buvy = wuky != cega;
	assign  xuqu = !(!vonu);
	assign  baxe = !abon ? !cyvu : 'z;
	assign  aras = !abon ? !bore : 'z;
	assign  agag = !abon ? !buvy : 'z;
	assign  abem = !abon ? !xuqu : 'z;
	assign  dyso = !abon ? !0 : 'z;
	assign  fufo = !ff40_d2;
	assign   gejy = (!xuso && fufo) || (ff40_d2 && wago);
	assign  famu = !abon ? !gejy : 'z;
	assign d[1] = xele;
	assign d[2] = ypon;
	assign d[3] = xuvo;
	assign d[4] = zysa;
	assign d[5] = yweg;
	assign d[6] = xabu;
	assign d[7] = ytux;
	assign d[0] = yfap;
	assign nma[5]  = fugy;
	assign nma[6]  = gavo;
	assign nma[7]  = wyga;
	assign nma[8]  = wune;
	assign nma[9]  = gotu;
	assign nma[10] = gegu;
	assign nma[11] = xehe;
	assign nma[1]  = baxe;
	assign nma[2]  = aras;
	assign nma[3]  = agag;
	assign nma[0]  = abem;
	assign nma[12] = dyso;
	assign nma[4]  = famu;
	assign spr_match = gese;

	logic xyva, xota, xyfy, wuvu, ales, abov, balu, wosu, bagy, wojo, ceno, byba;
	logic ceha, doba, care, bebu, dyty;
	dffr_bp dffr_wuvu(xota, nreset_video, !wuvu, wuvu);
	dffr_bp dffr_wosu(xyfy, nreset_video, !wuvu, wosu);
	dffr_bp dffr_ceno(xupy, abez,         besu,  ceno);
	dffr_bp dffr_catu(xupy, abez,         abov,  catu);
	dffr_bp dffr_byba(xupy, bagy,         feto,  byba);
	dffr_bp dffr_doba(clk2, bagy,         byba,  doba);
	assign  xyva = !clk1;
	assign  xota = !xyva;
	assign  xyfy = !xota;
	assign  ales = !xyvo;
	assign  abov = sela && ales;
	assign  balu = !anom;
	assign  xupy = !(!wuvu);
	assign  abez = !reset_video;
	assign  bagy = !balu;
	assign  wojo = !(!wosu || !wuvu);
	assign  xoce = !wosu;
	assign  xyso = !wojo;
	assign  ceha = !(!ceno);
	assign  buza = !ceno && nxymu;
	assign  care = xoce && ceha && spr_match;
	assign   bebu = doba || balu || !byba;
	assign  dyty = !care;
	assign  avap = !bebu;
	assign wuvu_nq = !wuvu;

	logic seba, toxe, tuly, tese, tepa, tyfo, tyno, saky, tytu, toma;
	logic vusa, tyso, tame, sycu, topu, raca, vywa, peby, weny, nybe;
	dffr_bp dffr_seba(clk4,  nxymu, vonu,  seba);
	dffr_bp dffr_toxe(toma,  seca,  !toxe, toxe);
	dffr_bp dffr_tuly(!toxe, seca,  !tuly, tuly);
	dffr_bp dffr_tese(!tuly, seca,  !tese, tese);
	dffr_bp dffr_tyfo(clk4,  '1,    toxe,  tyfo);
	assign  tepa = !nxymu;
	assign tyno = !(toxe && seba && vonu);
	assign  saky = !(tuly || vonu);
	assign  tytu = !toxe;
	assign   vusa = !tyfo || tyno;
	assign   tyso = saky || tepa;
	assign  tuvo = !(tepa || tuly || tese);
	assign tame = !(tese && toxe);
	assign  sycu = !(tytu || tepa || tyfo);
	assign tacu = !(tytu && tyfo);
	assign  wuty = !vusa;
	assign  texy = !tyso;
	assign  topu = tuly && sycu;
	assign  raca = vonu && sycu;
	assign  xefy = !wuty;
	assign  xono = nbaxo && texy;
	assign toma = !(clk4 && tame);
	assign  vywa = !topu;
	assign  peby = !raca;
	assign  weny = !vywa;
	assign  nybe = !peby;
	assign  xado = !weny;
	assign  puco = !nybe;
	assign tyfo_nq = !tyfo;

	logic baky, dezy, cake, bese, cuxy, bego, dybe;
	logic eden, cypy, cape, caxu, fycu, fone, ekud, elyg;
	logic gebu, womu, guna, foco, dewy, dezo, dogu, cugu, cupe, cuva;
	logic wyxo, xujo, gape, guve, caho, cemy, cato, cado, cecu, byby;
	logic gyfo, weka, gyvo, gusa, buka, dyhu, decu, bede, duke, buco;
	dffr_bp dffr_dezy(clk1,  nreset_video, dyty,  dezy);
	dffr_bp dffr_bese(cake,  azyb,         !bese, bese);
	dffr_bp dffr_cuxy(!bese, azyb,         !cuxy, cuxy);
	dffr_bp dffr_bego(!cuxy, azyb,         !bego, bego);
	dffr_bp dffr_dybe(!bego, azyb,         !dybe, dybe);
	assign  baky = cuxy && dybe;
	assign   cake = baky || dezy;
	assign  eden = !bese;
	assign  cypy = !cuxy;
	assign  cape = !bego;
	assign  caxu = !dybe;
	assign  fycu = !eden;
	assign  fone = !cypy;
	assign  ekud = !cape;
	assign  elyg = !caxu;
	assign gebu = !(eden && fone && cape && caxu);
	assign womu = !(eden && fone && ekud && caxu);
	assign guna = !(fycu && fone && ekud && caxu);
	assign foco = !(fycu && fone && cape && caxu);
	assign dewy = !(eden && cypy && cape && elyg);
	assign dezo = !(eden && cypy && cape && caxu);
	assign dogu = !(fycu && cypy && cape && elyg);
	assign cugu = !(fycu && cypy && ekud && caxu);
	assign cupe = !(eden && cypy && ekud && caxu);
	assign cuva = !(fycu && cypy && cape && caxu);
	assign   wyxo = dyty || gebu;
	assign   xujo = dyty || womu;
	assign   gape = dyty || guna;
	assign   guve = dyty || foco;
	assign   caho = dyty || dewy;
	assign   cemy = dyty || dezo;
	assign   cato = dyty || dogu;
	assign   cado = dyty || cugu;
	assign   cecu = dyty || cupe;
	assign   byby = dyty || cuva;
	assign  gyfo = !wyxo;
	assign  weka = !xujo;
	assign  gyvo = !gape;
	assign  gusa = !guve;
	assign  buka = !caho;
	assign  dyhu = !cemy;
	assign  decu = !cato;
	assign  bede = !cado;
	assign  duke = !cecu;
	assign  buco = !byby;
	assign  cacu = !gyfo;
	assign  buzy = !gyfo;
	assign  fuke = !gyfo;
	assign  zape = !weka;
	assign  wuse = !weka;
	assign  zuru = !weka;
	assign  fefo = !gyvo;
	assign  gecy = !gyvo;
	assign  wabe = !gyvo;
	assign  feka = !gusa;
	assign  xyha = !gusa;
	assign  yfag = !gusa;
	assign  cexu = !buka;
	assign  akol = !buka;
	assign  bymy = !buka;
	assign  fuxu = !dyhu;
	assign  enob = !dyhu;
	assign  geny = !dyhu;
	assign  weme = !decu;
	assign  wufa = !decu;
	assign  faka = !decu;
	assign  cyla = !bede;
	assign  dymo = !bede;
	assign  bucy = !bede;
	assign  wofo = !duke;
	assign  wylu = !duke;
	assign  ewot = !duke;
	assign  asys = !buco;
	assign  ahof = !buco;
	assign  byvy = !buco;

endmodule
