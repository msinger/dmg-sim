`default_nettype none

module sprite_x_matchers(
		inout tri logic [7:0] d,
		input logic     [7:0] oam_a_nd, nh,

		input logic clk3, oam_a_cpu_nrd,
		input logic cota, dyna, fuxu, wupa, yfag, gafy, gecy, asys, doku, zape, xaho, wunu, wofo,
		input logic wuzo, cexu, dosy, weme, ejad, cyla, cacu, gamy,

		output logic ngomo, nbaxo, nyzos, ndepo, xeba, zako, ywos, zure, daje, cyco, cyvy, ewam,
		output logic ywap, ydot, ykok, ynaz, dama, feha, ytub, ylev, cogy, fyma, cehu, ekes
	);

	logic wyno, cyra, zuve, eced, xyky, yrum, ysex, yvel;
	logic xega, gomo, baxo, yzos, depo, ylor, zyty, zyve, zezy;
	logic cose, arop, xatu, bady, zago, zocy, ypur, yvok;
	logic xaca, xagu, xepu, xygu, xuna, deve, zeha, fyra;
	logic welo, xuny, wote, xako, xepe, ylah, zola, zulu;
	logic woju, yfun, wyza, ypuk, zogy, zeba, zaha, zoky;
	logic xomy, wuha, wyna, weco, xoly, xyba, xabe, xeka;
	logic yvap, xeny, xavu, xeva, yhok, ycah, ydaj, yvuz;
	logic fazu, faxe, exuk, fede, eraz, epum, erol, ehyn;
	logic ejot, esaj, ducu, ewud, duse, dagu, dyze, deso;
	logic dake, ceso, dyfu, cusy, dany, duko, desu, dazo;
	logic cola, boba, colu, bahu, edym, emyb, ebef, ewok;
	logic zoly, zogo, zecu, zesa, ycol, yrac, ymem, yvag;
	logic zare, zemu, zygo, zuzy, xosu, zuvu, xuco, zulo;
	logic ybed, zala, wyde, xepa, wedu, ygaj, zyjo, xury;
	logic zyku, zypu, xaha, zefe, xeju, zate, zaku, ybox;
	logic ezuf, enad, ebow, fyca, gavy, gypu, gady, gaza;
	logic duze, daga, dawu, ejaw, goho, gasu, gabu, gafe;
	logic ypod, yrop, ynep, yzof, xuvy, xere, xuzo, xexa;
	logic zywu, zuza, zejo, zeda, ymam, ytyp, yfop, yvac;
	logic cywe, dyby, dury, cuvy, fusa, faxa, fozy, fesy;
	logic bazy, cyle, ceva, bumy, guzo, gola, geve, gude;
	logic duhy, ejuf, enor, depy, foka, fyty, fuby, goxu;
	logic ceko, dety, dozo, cony, fuzu, feso, foky, fyva;

	dlatch_a latch_gomo(!xega, wyno, gomo);
	dlatch_a latch_baxo(!xega, cyra, baxo);
	dlatch_a latch_yzos(!xega, zuve, yzos);
	dlatch_a latch_depo(!xega, eced, depo);
	dlatch_a latch_ylor(!xega, xyky, ylor);
	dlatch_a latch_zyty(!xega, yrum, zyty);
	dlatch_a latch_zyve(!xega, ysex, zyve);
	dlatch_a latch_zezy(!xega, yvel, zezy);
	dlatch_b latch_wyno(clk3, oam_a_nd[4], wyno);
	dlatch_b latch_cyra(clk3, oam_a_nd[5], cyra);
	dlatch_b latch_zuve(clk3, oam_a_nd[6], zuve);
	dlatch_b latch_eced(clk3, oam_a_nd[7], eced);
	dlatch_b latch_xyky(clk3, oam_a_nd[0], xyky);
	dlatch_b latch_yrum(clk3, oam_a_nd[1], yrum);
	dlatch_b latch_ysex(clk3, oam_a_nd[2], ysex);
	dlatch_b latch_yvel(clk3, oam_a_nd[3], yvel);
	drlatch latch_welo(!fuxu, dyna, cose, welo);
	drlatch latch_xuny(!fuxu, dyna, arop, xuny);
	drlatch latch_wote(!fuxu, dyna, xatu, wote);
	drlatch latch_xako(!fuxu, dyna, bady, xako);
	drlatch latch_xepe(!fuxu, dyna, zago, xepe);
	drlatch latch_ylah(!fuxu, dyna, zocy, ylah);
	drlatch latch_zola(!fuxu, dyna, ypur, zola);
	drlatch latch_zulu(!fuxu, dyna, yvok, zulu);
	drlatch latch_xomy(!yfag, wupa, cose, xomy);
	drlatch latch_wuha(!yfag, wupa, arop, wuha);
	drlatch latch_wyna(!yfag, wupa, xatu, wyna);
	drlatch latch_weco(!yfag, wupa, bady, weco);
	drlatch latch_xoly(!yfag, wupa, zago, xoly);
	drlatch latch_xyba(!yfag, wupa, zocy, xyba);
	drlatch latch_xabe(!yfag, wupa, ypur, xabe);
	drlatch latch_xeka(!yfag, wupa, yvok, xeka);
	drlatch latch_fazu(!gecy, gafy, cose, fazu);
	drlatch latch_faxe(!gecy, gafy, arop, faxe);
	drlatch latch_exuk(!gecy, gafy, xatu, exuk);
	drlatch latch_fede(!gecy, gafy, bady, fede);
	drlatch latch_eraz(!gecy, gafy, zago, eraz);
	drlatch latch_epum(!gecy, gafy, zocy, epum);
	drlatch latch_erol(!gecy, gafy, ypur, erol);
	drlatch latch_ehyn(!gecy, gafy, yvok, ehyn);
	drlatch latch_dake(!asys, doku, cose, dake);
	drlatch latch_ceso(!asys, doku, arop, ceso);
	drlatch latch_dyfu(!asys, doku, xatu, dyfu);
	drlatch latch_cusy(!asys, doku, bady, cusy);
	drlatch latch_dany(!asys, doku, zago, dany);
	drlatch latch_duko(!asys, doku, zocy, duko);
	drlatch latch_desu(!asys, doku, ypur, desu);
	drlatch latch_dazo(!asys, doku, yvok, dazo);
	drlatch latch_zecu(!zape, xaho, cose, zecu);
	drlatch latch_zogo(!zape, xaho, arop, zogo);
	drlatch latch_zoly(!zape, xaho, xatu, zoly);
	drlatch latch_zesa(!zape, xaho, bady, zesa);
	drlatch latch_ycol(!zape, xaho, zago, ycol);
	drlatch latch_yrac(!zape, xaho, zocy, yrac);
	drlatch latch_ymem(!zape, xaho, ypur, ymem);
	drlatch latch_yvag(!zape, xaho, yvok, yvag);
	drlatch latch_ybed(!wofo, wunu, cose, ybed);
	drlatch latch_zala(!wofo, wunu, arop, zala);
	drlatch latch_wyde(!wofo, wunu, xatu, wyde);
	drlatch latch_xepa(!wofo, wunu, bady, xepa);
	drlatch latch_wedu(!wofo, wunu, zago, wedu);
	drlatch latch_ygaj(!wofo, wunu, zocy, ygaj);
	drlatch latch_zyjo(!wofo, wunu, ypur, zyjo);
	drlatch latch_xury(!wofo, wunu, yvok, xury);
	drlatch latch_ezuf(!cexu, wuzo, cose, ezuf);
	drlatch latch_enad(!cexu, wuzo, arop, enad);
	drlatch latch_ebow(!cexu, wuzo, xatu, ebow);
	drlatch latch_fyca(!cexu, wuzo, bady, fyca);
	drlatch latch_gavy(!cexu, wuzo, zago, gavy);
	drlatch latch_gypu(!cexu, wuzo, zocy, gypu);
	drlatch latch_gady(!cexu, wuzo, ypur, gady);
	drlatch latch_gaza(!cexu, wuzo, yvok, gaza);
	drlatch latch_ypod(!weme, dosy, cose, ypod);
	drlatch latch_yrop(!weme, dosy, arop, yrop);
	drlatch latch_ynep(!weme, dosy, xatu, ynep);
	drlatch latch_yzof(!weme, dosy, bady, yzof);
	drlatch latch_xuvy(!weme, dosy, zago, xuvy);
	drlatch latch_xere(!weme, dosy, zocy, xere);
	drlatch latch_xuzo(!weme, dosy, ypur, xuzo);
	drlatch latch_xexa(!weme, dosy, yvok, xexa);
	drlatch latch_cywe(!cyla, ejad, cose, cywe);
	drlatch latch_dyby(!cyla, ejad, arop, dyby);
	drlatch latch_dury(!cyla, ejad, xatu, dury);
	drlatch latch_cuvy(!cyla, ejad, bady, cuvy);
	drlatch latch_fusa(!cyla, ejad, zago, fusa);
	drlatch latch_faxa(!cyla, ejad, zocy, faxa);
	drlatch latch_fozy(!cyla, ejad, ypur, fozy);
	drlatch latch_fesy(!cyla, ejad, yvok, fesy);
	drlatch latch_duhy(!cacu, gamy, cose, duhy);
	drlatch latch_ejuf(!cacu, gamy, arop, ejuf);
	drlatch latch_enor(!cacu, gamy, xatu, enor);
	drlatch latch_depy(!cacu, gamy, bady, depy);
	drlatch latch_foka(!cacu, gamy, zago, foka);
	drlatch latch_fyty(!cacu, gamy, zocy, fyty);
	drlatch latch_fuby(!cacu, gamy, ypur, fuby);
	drlatch latch_goxu(!cacu, gamy, yvok, goxu);
	assign #T_INV  xega = !cota;
	assign #T_INV  cose = !(!gomo);
	assign #T_INV  arop = !(!baxo);
	assign #T_INV  xatu = !(!yzos);
	assign #T_INV  bady = !(!depo);
	assign #T_INV  zago = !(!ylor);
	assign #T_INV  zocy = !(!zyty);
	assign #T_INV  ypur = !(!zyve);
	assign #T_INV  yvok = !(!zezy);
	assign #T_TRIB xaca = !oam_a_cpu_nrd ? !xyky : 'z;
	assign #T_TRIB xagu = !oam_a_cpu_nrd ? !yrum : 'z;
	assign #T_TRIB xepu = !oam_a_cpu_nrd ? !ysex : 'z;
	assign #T_TRIB xygu = !oam_a_cpu_nrd ? !yvel : 'z;
	assign #T_TRIB xuna = !oam_a_cpu_nrd ? !wyno : 'z;
	assign #T_TRIB deve = !oam_a_cpu_nrd ? !cyra : 'z;
	assign #T_TRIB zeha = !oam_a_cpu_nrd ? !zuve : 'z;
	assign #T_TRIB fyra = !oam_a_cpu_nrd ? !eced : 'z;
	assign #T_XOR  woju = welo != nh[4];
	assign #T_XOR  yfun = xuny != nh[5];
	assign #T_XOR  wyza = wote != nh[6];
	assign #T_XOR  ypuk = xako != nh[7];
	assign #T_XOR  zogy = xepe != nh[0];
	assign #T_XOR  zeba = ylah != nh[1];
	assign #T_XOR  zaha = zola != nh[2];
	assign #T_XOR  zoky = zulu != nh[3];
	assign #T_NOR  xeba = !(woju || yfun || wyza || ypuk);
	assign #T_NOR  zako = !(zogy || zeba || zaha || zoky);
	assign #T_XOR  yvap = xomy != nh[4];
	assign #T_XOR  xeny = wuha != nh[5];
	assign #T_XOR  xavu = wyna != nh[6];
	assign #T_XOR  xeva = weco != nh[7];
	assign #T_XOR  yhok = xoly != nh[0];
	assign #T_XOR  ycah = xyba != nh[1];
	assign #T_XOR  ydaj = xabe != nh[2];
	assign #T_XOR  yvuz = xeka != nh[3];
	assign #T_NOR  ywos = !(yvap || xeny || xavu || xeva);
	assign #T_NOR  zure = !(yhok || ycah || ydaj || yvuz);
	assign #T_XOR  ejot = fazu != nh[4];
	assign #T_XOR  esaj = faxe != nh[5];
	assign #T_XOR  ducu = exuk != nh[6];
	assign #T_XOR  ewud = fede != nh[7];
	assign #T_XOR  duse = eraz != nh[0];
	assign #T_XOR  dagu = epum != nh[1];
	assign #T_XOR  dyze = erol != nh[2];
	assign #T_XOR  deso = ehyn != nh[3];
	assign #T_NOR  daje = !(ejot || esaj || ducu || ewud);
	assign #T_NOR  cyco = !(duse || dagu || dyze || deso);
	assign #T_XOR  cola = dake != nh[4];
	assign #T_XOR  boba = ceso != nh[5];
	assign #T_XOR  colu = dyfu != nh[6];
	assign #T_XOR  bahu = cusy != nh[7];
	assign #T_XOR  edym = dany != nh[0];
	assign #T_XOR  emyb = duko != nh[1];
	assign #T_XOR  ebef = desu != nh[2];
	assign #T_XOR  ewok = dazo != nh[3];
	assign #T_NOR  cyvy = !(cola || boba || colu || bahu);
	assign #T_NOR  ewam = !(edym || emyb || ebef || ewok);
	assign #T_XOR  zare = zoly != nh[6];
	assign #T_XOR  zemu = zogo != nh[5];
	assign #T_XOR  zygo = zecu != nh[4];
	assign #T_XOR  zuzy = zesa != nh[7];
	assign #T_XOR  xosu = ycol != nh[0];
	assign #T_XOR  zuvu = yrac != nh[1];
	assign #T_XOR  xuco = ymem != nh[2];
	assign #T_XOR  zulo = yvag != nh[3];
	assign #T_NOR  ywap = !(zare || zemu || zygo || zuzy);
	assign #T_NOR  ydot = !(xosu || zuvu || xuco || zulo);
	assign #T_XOR  zyku = ybed != nh[4];
	assign #T_XOR  zypu = zala != nh[5];
	assign #T_XOR  xaha = wyde != nh[6];
	assign #T_XOR  zefe = xepa != nh[7];
	assign #T_XOR  xeju = wedu != nh[0];
	assign #T_XOR  zate = ygaj != nh[1];
	assign #T_XOR  zaku = zyjo != nh[2];
	assign #T_XOR  ybox = xury != nh[3];
	assign #T_NOR  ykok = !(zyku || zypu || xaha || zefe);
	assign #T_NOR  ynaz = !(xeju || zate || zaku || ybox);
	assign #T_XOR  duze = ezuf != nh[4];
	assign #T_XOR  daga = enad != nh[5];
	assign #T_XOR  dawu = ebow != nh[6];
	assign #T_XOR  ejaw = fyca != nh[7];
	assign #T_XOR  goho = gavy != nh[0];
	assign #T_XOR  gasu = gypu != nh[1];
	assign #T_XOR  gabu = gady != nh[2];
	assign #T_XOR  gafe = gaza != nh[3];
	assign #T_NOR  dama = !(duze || daga || dawu || ejaw);
	assign #T_NOR  feha = !(goho || gasu || gabu || gafe);
	assign #T_XOR  zywu = ypod != nh[4];
	assign #T_XOR  zuza = yrop != nh[5];
	assign #T_XOR  zejo = ynep != nh[6];
	assign #T_XOR  zeda = yzof != nh[7];
	assign #T_XOR  ymam = xuvy != nh[0];
	assign #T_XOR  ytyp = xere != nh[1];
	assign #T_XOR  yfop = xuzo != nh[2];
	assign #T_XOR  yvac = xexa != nh[3];
	assign #T_NOR  ytub = !(zywu || zuza || zejo || zeda);
	assign #T_NOR  ylev = !(ymam || ytyp || yfop || yvac);
	assign #T_XOR  bazy = cywe != nh[4];
	assign #T_XOR  cyle = dyby != nh[5];
	assign #T_XOR  ceva = dury != nh[6];
	assign #T_XOR  bumy = cuvy != nh[7];
	assign #T_XOR  guzo = fusa != nh[0];
	assign #T_XOR  gola = faxa != nh[1];
	assign #T_XOR  geve = fozy != nh[2];
	assign #T_XOR  gude = fesy != nh[3];
	assign #T_NOR  cogy = !(bazy || cyle || ceva || bumy);
	assign #T_NOR  fyma = !(guzo || gola || geve || gude);
	assign #T_XOR  ceko = duhy != nh[4];
	assign #T_XOR  dety = ejuf != nh[5];
	assign #T_XOR  dozo = enor != nh[6];
	assign #T_XOR  cony = depy != nh[7];
	assign #T_XOR  fuzu = foka != nh[0];
	assign #T_XOR  feso = fyty != nh[1];
	assign #T_XOR  foky = fuby != nh[2];
	assign #T_XOR  fyva = goxu != nh[3];
	assign #T_NOR  cehu = !(ceko || dety || dozo || cony);
	assign #T_NOR  ekes = !(fuzu || feso || foky || fyva);
	assign ngomo = !gomo;
	assign nbaxo = !baxo;
	assign nyzos = !yzos;
	assign ndepo = !depo;
	assign d[0] = xaca;
	assign d[1] = xagu;
	assign d[2] = xepu;
	assign d[3] = xygu;
	assign d[4] = xuna;
	assign d[5] = deve;
	assign d[6] = zeha;
	assign d[7] = fyra;

endmodule
