`default_nettype none

module sprite_pixel_shifter(
		input  logic [7:0] md,
		output logic [7:0] spr_pix_a, spr_pix_b,

		input logic clkpipe, xono, xado, puco,
		input logic roby, lyku, lesy, lota, tyta, tyco, xovu, soka
	);

	logic pobe, pacy, pono, pugu, pute, puly, pelo, pawe;
	logic pudu, ramu, mytu, mofo, pefo, rewo, peba, roka;
	logic lubo, solo, lumo, lase, loza, rata, nuca, sybo;
	logic lufy, mame, rehu, rano, majo, myxa, lyde, lela;
	logic mofy, mezu, pyzu, pabe, mada, myto, ruca, rusy;
	logic sele, saja, suny, suto, rydu, sega, rama, semo;
	logic voby, wery, wura, wyco, selu, wamy, sery, sulu;
	logic waxo, tyga, xato, vexu, xexu, vaby, xole, vume;
	logic tula, teso, xyve, vune, taby, tapo, tupe, tuxa;
	dlatch_a latch_pudu(!xado, pobe, pudu);
	dlatch_a latch_ramu(!puco, pobe, ramu);
	dlatch_a latch_mytu(!puco, pono, mytu);
	dlatch_a latch_mofo(!xado, pono, mofo);
	dlatch_a latch_pefo(!puco, pute, pefo);
	dlatch_a latch_rewo(!xado, pute, rewo);
	dlatch_a latch_peba(!xado, pelo, peba);
	dlatch_a latch_roka(!puco, pelo, roka);
	dlatch_a latch_sele(!puco, pacy, sele);
	dlatch_a latch_saja(!xado, pacy, saja);
	dlatch_a latch_suny(!xado, pugu, suny);
	dlatch_a latch_suto(!puco, pugu, suto);
	dlatch_a latch_rydu(!puco, puly, rydu);
	dlatch_a latch_sega(!xado, puly, sega);
	dlatch_a latch_rama(!puco, pawe, rama);
	dlatch_a latch_semo(!xado, pawe, semo);
	assign  pobe = xono ? md[4] : md[3];
	assign  pacy = xono ? md[3] : md[4];
	assign  pono = xono ? md[5] : md[2];
	assign  pugu = xono ? md[2] : md[5];
	assign  pute = xono ? md[7] : md[0];
	assign  puly = xono ? md[0] : md[7];
	assign  pelo = xono ? md[6] : md[1];
	assign  pawe = xono ? md[1] : md[6];
	assign  lubo = !pudu;
	assign  solo = !ramu;
	assign  lumo = !mytu;
	assign  lase = !mofo;
	assign  loza = !pefo;
	assign  rata = !rewo;
	assign  nuca = !peba;
	assign  sybo = !roka;
	assign lufy = !(lubo && roby);
	assign mame = !(pudu && roby);
	assign rehu = !(solo && roby);
	assign rano = !(ramu && roby);
	assign majo = !(lumo && lyku);
	assign myxa = !(mytu && lyku);
	assign lyde = !(lase && lyku);
	assign lela = !(mofo && lyku);
	assign mofy = !(loza && lesy);
	assign mezu = !(pefo && lesy);
	assign pyzu = !(rata && lesy);
	assign pabe = !(rewo && lesy);
	assign mada = !(nuca && lota);
	assign myto = !(peba && lota);
	assign ruca = !(sybo && lota);
	assign rusy = !(roka && lota);
	assign  voby = !sele;
	assign  wery = !saja;
	assign  wura = !suny;
	assign  wyco = !suto;
	assign  selu = !rydu;
	assign  wamy = !sega;
	assign  sery = !rama;
	assign  sulu = !semo;
	assign waxo = !(voby && tyta);
	assign tyga = !(sele && tyta);
	assign xato = !(wery && tyta);
	assign vexu = !(saja && tyta);
	assign xexu = !(wura && tyco);
	assign vaby = !(suny && tyco);
	assign xole = !(wyco && tyco);
	assign vume = !(suto && tyco);
	assign tula = !(selu && xovu);
	assign teso = !(rydu && xovu);
	assign xyve = !(wamy && xovu);
	assign vune = !(sega && xovu);
	assign taby = !(sery && soka);
	assign tapo = !(rama && soka);
	assign tupe = !(sulu && soka);
	assign tuxa = !(semo && soka);
	assign  pobe = xono ? md[4] : md[3];
	assign  pacy = xono ? md[3] : md[4];
	assign  pono = xono ? md[5] : md[2];
	assign  pugu = xono ? md[2] : md[5];
	assign  pute = xono ? md[7] : md[0];
	assign  puly = xono ? md[0] : md[7];
	assign  pelo = xono ? md[6] : md[1];
	assign  pawe = xono ? md[1] : md[6];
	assign  lubo = !pudu;
	assign  solo = !ramu;
	assign  lumo = !mytu;
	assign  lase = !mofo;
	assign  loza = !pefo;
	assign  rata = !rewo;
	assign  nuca = !peba;
	assign  sybo = !roka;
	assign lufy = !(lubo && roby);
	assign mame = !(pudu && roby);
	assign rehu = !(solo && roby);
	assign rano = !(ramu && roby);
	assign majo = !(lumo && lyku);
	assign myxa = !(mytu && lyku);
	assign lyde = !(lase && lyku);
	assign lela = !(mofo && lyku);
	assign mofy = !(loza && lesy);
	assign mezu = !(pefo && lesy);
	assign pyzu = !(rata && lesy);
	assign pabe = !(rewo && lesy);
	assign mada = !(nuca && lota);
	assign myto = !(peba && lota);
	assign ruca = !(sybo && lota);
	assign rusy = !(roka && lota);
	assign  voby = !sele;
	assign  wery = !saja;
	assign  wura = !suny;
	assign  wyco = !suto;
	assign  selu = !rydu;
	assign  wamy = !sega;
	assign  sery = !sery;
	assign  sulu = !semo;
	assign waxo = !(voby && tyta);
	assign tyga = !(sele && tyta);
	assign xato = !(wery && tyta);
	assign vexu = !(saja && tyta);
	assign xexu = !(wura && tyco);
	assign vaby = !(suny && tyco);
	assign xole = !(wyco && tyco);
	assign vume = !(suto && tyco);
	assign tula = !(selu && xovu);
	assign teso = !(rydu && xovu);
	assign xyve = !(wamy && xovu);
	assign vune = !(sega && xovu);
	assign taby = !(sery && soka);
	assign tapo = !(rama && soka);
	assign tupe = !(sulu && soka);
	assign tuxa = !(semo && soka);

	logic nuro, maso, lefe, lesu, wyho, wora, vafo, wufy;
	logic nylu, pefu, naty, pyjo, vare, weba, vanu, vupy;
	dffsr dffsr_nuro(clkpipe, pabe, pyzu, '0,   nuro);
	dffsr dffsr_maso(clkpipe, myto, mada, nuro, maso);
	dffsr dffsr_lefe(clkpipe, lela, lyde, maso, lefe);
	dffsr dffsr_lesu(clkpipe, mame, lufy, lefe, lesu);
	dffsr dffsr_wyho(clkpipe, vexu, xato, lesu, wyho);
	dffsr dffsr_wora(clkpipe, vaby, xexu, wyho, wora);
	dffsr dffsr_vafo(clkpipe, tuxa, tupe, wora, vafo);
	dffsr dffsr_wufy(clkpipe, vune, xyve, vafo, wufy);
	dffsr dffsr_nylu(clkpipe, mezu, mofy, '0,   nylu);
	dffsr dffsr_pefu(clkpipe, rusy, ruca, nylu, pefu);
	dffsr dffsr_naty(clkpipe, myxa, majo, pefu, naty);
	dffsr dffsr_pyjo(clkpipe, rano, rehu, naty, pyjo);
	dffsr dffsr_vare(clkpipe, tyga, waxo, pyjo, vare);
	dffsr dffsr_weba(clkpipe, vume, xole, vare, weba);
	dffsr dffsr_vanu(clkpipe, tapo, taby, weba, vanu);
	dffsr dffsr_vupy(clkpipe, teso, tula, vanu, vupy);
	assign spr_pix_b[0] = nuro;
	assign spr_pix_b[1] = maso;
	assign spr_pix_b[2] = lefe;
	assign spr_pix_b[3] = lesu;
	assign spr_pix_b[4] = wyho;
	assign spr_pix_b[5] = wora;
	assign spr_pix_b[6] = vafo;
	assign spr_pix_b[7] = wufy;
	assign spr_pix_a[0] = nylu;
	assign spr_pix_a[1] = pefu;
	assign spr_pix_a[2] = naty;
	assign spr_pix_a[3] = pyjo;
	assign spr_pix_a[4] = vare;
	assign spr_pix_a[5] = weba;
	assign spr_pix_a[6] = vanu;
	assign spr_pix_a[7] = vupy;

endmodule
