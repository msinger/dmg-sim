`default_nettype none

parameter time T_INV     = 2ns;
parameter time T_AND     = 4ns;
parameter time T_NAND    = 2ns;
parameter time T_OR      = 4ns;
parameter time T_NOR     = 2ns;
parameter time T_OA      = 6ns;
parameter time T_AO      = 6ns;
parameter time T_NAO     = 5ns;
parameter time T_MUX     = 6ns;
parameter time T_MUXI    = 6ns;
parameter time T_AOI     = 5ns;
parameter time T_XOR     = 5ns;
parameter time T_XNOR    = 5ns;
parameter time T_ADD     = 6ns;
parameter time T_TRI     = 2ns;
parameter time T_SRL     = 4ns;
parameter time T_DL      = 4ns;
parameter time T_DFF     = 8ns;
parameter time T_DFFR_A  = 8ns;
parameter time T_DFFR_B  = 8ns;
parameter time T_DFFR_BP = 8ns;
parameter time T_DFFR_C  = 8ns;
parameter time T_DFFSR   = 8ns;
parameter time T_TFFD    = 8ns;
