`default_nettype none

parameter time T_INV   = 2ns;
parameter time T_AND   = 4ns;
parameter time T_NAND  = 2ns;
parameter time T_OR    = 4ns;
parameter time T_NOR   = 2ns;
parameter time T_OA    = 6ns;
parameter time T_AO    = 6ns;
parameter time T_NAO   = 5ns;
parameter time T_MUX   = 6ns;
parameter time T_MUXI  = 6ns;
parameter time T_AOI   = 5ns;
parameter time T_XOR   = 5ns;
parameter time T_ADD   = 6ns;
parameter time T_TRI   = 2ns;
parameter time T_DFFSR = 8ns;
parameter time T_DFFR  = 8ns;
parameter time T_DFF   = 8ns;
parameter time T_LATCH = 4ns;
parameter time T_COUNT = 8ns;
